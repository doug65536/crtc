module crt (clk, reset, cs, we, addr, data, irq, vs, hs, ven, clksel, pixaddr);

input clk;
input reset;
input cs;
input we;
output irq;
output vs;
output hs;
output ven;
input [3:0] addr;
input [15:0] data;
output [2:0] clksel;
output [31:0] pixaddr;

wire vdd = 1'b1;
wire gnd = 1'b0;

	INVX8 INVX8_1 ( .A(reset), .Y(_abc_3927_n365) );
	XNOR2X1 XNOR2X1_1 ( .A(currentrow_10_), .B(reg_ve_value_10_), .Y(_abc_3927_n366) );
	XNOR2X1 XNOR2X1_2 ( .A(currentrow_11_), .B(reg_ve_value_11_), .Y(_abc_3927_n367) );
	NAND2X1 NAND2X1_1 ( .A(_abc_3927_n366), .B(_abc_3927_n367), .Y(_abc_3927_n368) );
	XNOR2X1 XNOR2X1_3 ( .A(currentrow_14_), .B(reg_ve_value_14_), .Y(_abc_3927_n369) );
	INVX1 INVX1_1 ( .A(_abc_3927_n369), .Y(_abc_3927_n370) );
	XOR2X1 XOR2X1_1 ( .A(currentrow_15_), .B(reg_ve_value_15_), .Y(_abc_3927_n371) );
	NOR2X1 NOR2X1_1 ( .A(_abc_3927_n371), .B(_abc_3927_n370), .Y(_abc_3927_n372) );
	INVX1 INVX1_2 ( .A(_abc_3927_n372), .Y(_abc_3927_n373) );
	NOR2X1 NOR2X1_2 ( .A(_abc_3927_n368), .B(_abc_3927_n373), .Y(_abc_3927_n374) );
	XNOR2X1 XNOR2X1_4 ( .A(currentrow_1_), .B(reg_ve_value_1_), .Y(_abc_3927_n375) );
	XNOR2X1 XNOR2X1_5 ( .A(currentrow_0_), .B(reg_ve_value_0_), .Y(_abc_3927_n376) );
	NAND2X1 NAND2X1_2 ( .A(_abc_3927_n375), .B(_abc_3927_n376), .Y(_abc_3927_n377) );
	XOR2X1 XOR2X1_2 ( .A(currentrow_4_), .B(reg_ve_value_4_), .Y(_abc_3927_n378) );
	XOR2X1 XOR2X1_3 ( .A(currentrow_5_), .B(reg_ve_value_5_), .Y(_abc_3927_n379) );
	NOR2X1 NOR2X1_3 ( .A(_abc_3927_n378), .B(_abc_3927_n379), .Y(_abc_3927_n380) );
	INVX1 INVX1_3 ( .A(_abc_3927_n380), .Y(_abc_3927_n381) );
	NOR2X1 NOR2X1_4 ( .A(_abc_3927_n377), .B(_abc_3927_n381), .Y(_abc_3927_n382) );
	NAND2X1 NAND2X1_3 ( .A(_abc_3927_n382), .B(_abc_3927_n374), .Y(_abc_3927_n383) );
	XNOR2X1 XNOR2X1_6 ( .A(currentrow_8_), .B(reg_ve_value_8_), .Y(_abc_3927_n384) );
	XNOR2X1 XNOR2X1_7 ( .A(currentrow_9_), .B(reg_ve_value_9_), .Y(_abc_3927_n385) );
	NAND2X1 NAND2X1_4 ( .A(_abc_3927_n384), .B(_abc_3927_n385), .Y(_abc_3927_n386) );
	XOR2X1 XOR2X1_4 ( .A(currentrow_13_), .B(reg_ve_value_13_), .Y(_abc_3927_n387) );
	XOR2X1 XOR2X1_5 ( .A(currentrow_12_), .B(reg_ve_value_12_), .Y(_abc_3927_n388) );
	NOR2X1 NOR2X1_5 ( .A(_abc_3927_n387), .B(_abc_3927_n388), .Y(_abc_3927_n389) );
	INVX1 INVX1_4 ( .A(_abc_3927_n389), .Y(_abc_3927_n390) );
	NOR2X1 NOR2X1_6 ( .A(_abc_3927_n386), .B(_abc_3927_n390), .Y(_abc_3927_n391) );
	INVX1 INVX1_5 ( .A(_abc_3927_n391), .Y(_abc_3927_n392) );
	XNOR2X1 XNOR2X1_8 ( .A(currentrow_3_), .B(reg_ve_value_3_), .Y(_abc_3927_n393) );
	INVX1 INVX1_6 ( .A(_abc_3927_n393), .Y(_abc_3927_n394) );
	XOR2X1 XOR2X1_6 ( .A(currentrow_2_), .B(reg_ve_value_2_), .Y(_abc_3927_n395) );
	NOR2X1 NOR2X1_7 ( .A(_abc_3927_n395), .B(_abc_3927_n394), .Y(_abc_3927_n396) );
	XNOR2X1 XNOR2X1_9 ( .A(currentrow_7_), .B(reg_ve_value_7_), .Y(_abc_3927_n397) );
	INVX1 INVX1_7 ( .A(_abc_3927_n397), .Y(_abc_3927_n398) );
	XOR2X1 XOR2X1_7 ( .A(currentrow_6_), .B(reg_ve_value_6_), .Y(_abc_3927_n399) );
	NOR2X1 NOR2X1_8 ( .A(_abc_3927_n399), .B(_abc_3927_n398), .Y(_abc_3927_n400) );
	NAND2X1 NAND2X1_5 ( .A(_abc_3927_n396), .B(_abc_3927_n400), .Y(_abc_3927_n401) );
	NOR2X1 NOR2X1_9 ( .A(_abc_3927_n401), .B(_abc_3927_n392), .Y(_abc_3927_n402) );
	INVX1 INVX1_8 ( .A(_abc_3927_n402), .Y(_abc_3927_n403) );
	NOR2X1 NOR2X1_10 ( .A(_abc_3927_n383), .B(_abc_3927_n403), .Y(_abc_3927_n404) );
	INVX8 INVX8_2 ( .A(_abc_3927_n404), .Y(_abc_3927_n405) );
	INVX1 INVX1_9 ( .A(currentaddr_30_), .Y(_abc_3927_n406) );
	INVX2 INVX2_1 ( .A(currentaddr_28_), .Y(_abc_3927_n407) );
	INVX1 INVX1_10 ( .A(currentaddr_29_), .Y(_abc_3927_n408) );
	NOR2X1 NOR2X1_11 ( .A(_abc_3927_n407), .B(_abc_3927_n408), .Y(_abc_3927_n409) );
	INVX1 INVX1_11 ( .A(currentaddr_25_), .Y(_abc_3927_n410) );
	INVX1 INVX1_12 ( .A(currentaddr_24_), .Y(_abc_3927_n411) );
	NOR2X1 NOR2X1_12 ( .A(_abc_3927_n410), .B(_abc_3927_n411), .Y(_abc_3927_n412) );
	INVX1 INVX1_13 ( .A(currentaddr_27_), .Y(_abc_3927_n413) );
	INVX2 INVX2_2 ( .A(currentaddr_26_), .Y(_abc_3927_n414) );
	NOR2X1 NOR2X1_13 ( .A(_abc_3927_n413), .B(_abc_3927_n414), .Y(_abc_3927_n415) );
	NAND2X1 NAND2X1_6 ( .A(_abc_3927_n412), .B(_abc_3927_n415), .Y(_abc_3927_n416) );
	INVX1 INVX1_14 ( .A(_abc_3927_n416), .Y(_abc_3927_n417) );
	AND2X2 AND2X2_1 ( .A(_abc_3927_n417), .B(_abc_3927_n409), .Y(_abc_3927_n418) );
	INVX2 INVX2_3 ( .A(currentrow_15_), .Y(_abc_3927_n419) );
	NAND2X1 NAND2X1_7 ( .A(reg_vf_value_15_), .B(_abc_3927_n419), .Y(_abc_3927_n420) );
	OR2X2 OR2X2_1 ( .A(_abc_3927_n419), .B(reg_vf_value_15_), .Y(_abc_3927_n421) );
	AND2X2 AND2X2_2 ( .A(_abc_3927_n421), .B(_abc_3927_n420), .Y(_abc_3927_n422) );
	INVX2 INVX2_4 ( .A(currentrow_14_), .Y(_abc_3927_n423) );
	AND2X2 AND2X2_3 ( .A(_abc_3927_n423), .B(reg_vf_value_14_), .Y(_abc_3927_n424) );
	NOR2X1 NOR2X1_14 ( .A(reg_vf_value_14_), .B(_abc_3927_n423), .Y(_abc_3927_n425) );
	NOR2X1 NOR2X1_15 ( .A(_abc_3927_n425), .B(_abc_3927_n424), .Y(_abc_3927_n426_1) );
	NAND2X1 NAND2X1_8 ( .A(_abc_3927_n426_1), .B(_abc_3927_n422), .Y(_abc_3927_n427_1) );
	INVX2 INVX2_5 ( .A(currentrow_12_), .Y(_abc_3927_n428_1) );
	NOR2X1 NOR2X1_16 ( .A(reg_vf_value_12_), .B(_abc_3927_n428_1), .Y(_abc_3927_n429_1) );
	AND2X2 AND2X2_4 ( .A(_abc_3927_n428_1), .B(reg_vf_value_12_), .Y(_abc_3927_n430_1) );
	NOR2X1 NOR2X1_17 ( .A(_abc_3927_n429_1), .B(_abc_3927_n430_1), .Y(_abc_3927_n431_1) );
	INVX2 INVX2_6 ( .A(currentrow_13_), .Y(_abc_3927_n432_1) );
	NOR2X1 NOR2X1_18 ( .A(reg_vf_value_13_), .B(_abc_3927_n432_1), .Y(_abc_3927_n433_1) );
	AND2X2 AND2X2_5 ( .A(_abc_3927_n432_1), .B(reg_vf_value_13_), .Y(_abc_3927_n434_1) );
	NOR2X1 NOR2X1_19 ( .A(_abc_3927_n433_1), .B(_abc_3927_n434_1), .Y(_abc_3927_n435_1) );
	NAND2X1 NAND2X1_9 ( .A(_abc_3927_n431_1), .B(_abc_3927_n435_1), .Y(_abc_3927_n436_1) );
	OR2X2 OR2X2_2 ( .A(_abc_3927_n427_1), .B(_abc_3927_n436_1), .Y(_abc_3927_n437_1) );
	INVX2 INVX2_7 ( .A(currentrow_11_), .Y(_abc_3927_n438_1) );
	NAND2X1 NAND2X1_10 ( .A(reg_vf_value_11_), .B(_abc_3927_n438_1), .Y(_abc_3927_n439_1) );
	OR2X2 OR2X2_3 ( .A(_abc_3927_n438_1), .B(reg_vf_value_11_), .Y(_abc_3927_n440_1) );
	NAND2X1 NAND2X1_11 ( .A(_abc_3927_n439_1), .B(_abc_3927_n440_1), .Y(_abc_3927_n441) );
	XOR2X1 XOR2X1_8 ( .A(reg_vf_value_10_), .B(currentrow_10_), .Y(_abc_3927_n442) );
	NOR2X1 NOR2X1_20 ( .A(_abc_3927_n442), .B(_abc_3927_n441), .Y(_abc_3927_n443) );
	INVX1 INVX1_15 ( .A(reg_vf_value_8_), .Y(_abc_3927_n444) );
	NAND2X1 NAND2X1_12 ( .A(currentrow_8_), .B(_abc_3927_n444), .Y(_abc_3927_n445) );
	INVX2 INVX2_8 ( .A(currentrow_9_), .Y(_abc_3927_n446) );
	OR2X2 OR2X2_4 ( .A(_abc_3927_n446), .B(reg_vf_value_9_), .Y(_abc_3927_n447) );
	NAND2X1 NAND2X1_13 ( .A(_abc_3927_n445), .B(_abc_3927_n447), .Y(_abc_3927_n448) );
	NOR2X1 NOR2X1_21 ( .A(currentrow_8_), .B(_abc_3927_n444), .Y(_abc_3927_n449) );
	INVX1 INVX1_16 ( .A(_abc_3927_n449), .Y(_abc_3927_n450) );
	NAND2X1 NAND2X1_14 ( .A(reg_vf_value_9_), .B(_abc_3927_n446), .Y(_abc_3927_n451_1) );
	NAND2X1 NAND2X1_15 ( .A(_abc_3927_n451_1), .B(_abc_3927_n450), .Y(_abc_3927_n452_1) );
	NOR2X1 NOR2X1_22 ( .A(_abc_3927_n448), .B(_abc_3927_n452_1), .Y(_abc_3927_n453) );
	NAND2X1 NAND2X1_16 ( .A(_abc_3927_n443), .B(_abc_3927_n453), .Y(_abc_3927_n454) );
	OR2X2 OR2X2_5 ( .A(_abc_3927_n437_1), .B(_abc_3927_n454), .Y(_abc_3927_n455) );
	INVX2 INVX2_9 ( .A(currentrow_7_), .Y(_abc_3927_n456) );
	NAND2X1 NAND2X1_17 ( .A(reg_vf_value_7_), .B(_abc_3927_n456), .Y(_abc_3927_n457) );
	OR2X2 OR2X2_6 ( .A(_abc_3927_n456), .B(reg_vf_value_7_), .Y(_abc_3927_n458) );
	NAND2X1 NAND2X1_18 ( .A(_abc_3927_n457), .B(_abc_3927_n458), .Y(_abc_3927_n459) );
	XOR2X1 XOR2X1_9 ( .A(reg_vf_value_6_), .B(currentrow_6_), .Y(_abc_3927_n460) );
	NOR2X1 NOR2X1_23 ( .A(_abc_3927_n460), .B(_abc_3927_n459), .Y(_abc_3927_n461) );
	INVX2 INVX2_10 ( .A(currentrow_5_), .Y(_abc_3927_n462) );
	OR2X2 OR2X2_7 ( .A(_abc_3927_n462), .B(reg_vf_value_5_), .Y(_abc_3927_n463) );
	INVX1 INVX1_17 ( .A(currentrow_4_), .Y(_abc_3927_n464) );
	NAND2X1 NAND2X1_19 ( .A(reg_vf_value_4_), .B(_abc_3927_n464), .Y(_abc_3927_n465) );
	NAND2X1 NAND2X1_20 ( .A(_abc_3927_n465), .B(_abc_3927_n463), .Y(_abc_3927_n466) );
	OR2X2 OR2X2_8 ( .A(_abc_3927_n464), .B(reg_vf_value_4_), .Y(_abc_3927_n467) );
	NAND2X1 NAND2X1_21 ( .A(reg_vf_value_5_), .B(_abc_3927_n462), .Y(_abc_3927_n468) );
	NAND2X1 NAND2X1_22 ( .A(_abc_3927_n468), .B(_abc_3927_n467), .Y(_abc_3927_n469) );
	NOR2X1 NOR2X1_24 ( .A(_abc_3927_n466), .B(_abc_3927_n469), .Y(_abc_3927_n470) );
	AND2X2 AND2X2_6 ( .A(_abc_3927_n470), .B(_abc_3927_n461), .Y(_abc_3927_n471) );
	INVX2 INVX2_11 ( .A(currentrow_3_), .Y(_abc_3927_n472) );
	NAND2X1 NAND2X1_23 ( .A(reg_vf_value_3_), .B(_abc_3927_n472), .Y(_abc_3927_n473) );
	OR2X2 OR2X2_9 ( .A(_abc_3927_n472), .B(reg_vf_value_3_), .Y(_abc_3927_n474) );
	NAND2X1 NAND2X1_24 ( .A(_abc_3927_n473), .B(_abc_3927_n474), .Y(_abc_3927_n475) );
	XOR2X1 XOR2X1_10 ( .A(reg_vf_value_2_), .B(currentrow_2_), .Y(_abc_3927_n476) );
	NOR2X1 NOR2X1_25 ( .A(_abc_3927_n476), .B(_abc_3927_n475), .Y(_abc_3927_n477) );
	INVX1 INVX1_18 ( .A(currentrow_1_), .Y(_abc_3927_n478_1) );
	NAND2X1 NAND2X1_25 ( .A(reg_vf_value_1_), .B(_abc_3927_n478_1), .Y(_abc_3927_n479) );
	INVX2 INVX2_12 ( .A(currentrow_0_), .Y(_abc_3927_n480_1) );
	OR2X2 OR2X2_10 ( .A(_abc_3927_n480_1), .B(reg_vf_value_0_), .Y(_abc_3927_n481) );
	XNOR2X1 XNOR2X1_10 ( .A(reg_vf_value_1_), .B(currentrow_1_), .Y(_abc_3927_n482) );
	NAND2X1 NAND2X1_26 ( .A(_abc_3927_n481), .B(_abc_3927_n482), .Y(_abc_3927_n483_1) );
	NAND2X1 NAND2X1_27 ( .A(_abc_3927_n479), .B(_abc_3927_n483_1), .Y(_abc_3927_n484) );
	NAND2X1 NAND2X1_28 ( .A(_abc_3927_n477), .B(_abc_3927_n484), .Y(_abc_3927_n485) );
	INVX2 INVX2_13 ( .A(currentrow_2_), .Y(_abc_3927_n486_1) );
	AND2X2 AND2X2_7 ( .A(_abc_3927_n486_1), .B(reg_vf_value_2_), .Y(_abc_3927_n487) );
	NAND2X1 NAND2X1_29 ( .A(_abc_3927_n487), .B(_abc_3927_n474), .Y(_abc_3927_n488) );
	AND2X2 AND2X2_8 ( .A(_abc_3927_n488), .B(_abc_3927_n473), .Y(_abc_3927_n489_1) );
	NAND2X1 NAND2X1_30 ( .A(_abc_3927_n489_1), .B(_abc_3927_n485), .Y(_abc_3927_n490) );
	NAND2X1 NAND2X1_31 ( .A(_abc_3927_n471), .B(_abc_3927_n490), .Y(_abc_3927_n491) );
	INVX1 INVX1_19 ( .A(_abc_3927_n465), .Y(_abc_3927_n492) );
	NAND2X1 NAND2X1_32 ( .A(_abc_3927_n463), .B(_abc_3927_n492), .Y(_abc_3927_n493_1) );
	NAND2X1 NAND2X1_33 ( .A(_abc_3927_n468), .B(_abc_3927_n493_1), .Y(_abc_3927_n494) );
	AND2X2 AND2X2_9 ( .A(_abc_3927_n461), .B(_abc_3927_n494), .Y(_abc_3927_n495) );
	INVX1 INVX1_20 ( .A(currentrow_6_), .Y(_abc_3927_n496) );
	AND2X2 AND2X2_10 ( .A(_abc_3927_n496), .B(reg_vf_value_6_), .Y(_abc_3927_n497) );
	NAND2X1 NAND2X1_34 ( .A(_abc_3927_n497), .B(_abc_3927_n458), .Y(_abc_3927_n498) );
	NAND2X1 NAND2X1_35 ( .A(_abc_3927_n457), .B(_abc_3927_n498), .Y(_abc_3927_n499) );
	NOR2X1 NOR2X1_26 ( .A(_abc_3927_n499), .B(_abc_3927_n495), .Y(_abc_3927_n500) );
	AND2X2 AND2X2_11 ( .A(_abc_3927_n491), .B(_abc_3927_n500), .Y(_abc_3927_n501_1) );
	OR2X2 OR2X2_11 ( .A(_abc_3927_n501_1), .B(_abc_3927_n455), .Y(_abc_3927_n502) );
	NAND2X1 NAND2X1_36 ( .A(_abc_3927_n449), .B(_abc_3927_n447), .Y(_abc_3927_n503) );
	NAND2X1 NAND2X1_37 ( .A(_abc_3927_n451_1), .B(_abc_3927_n503), .Y(_abc_3927_n504_1) );
	AND2X2 AND2X2_12 ( .A(_abc_3927_n443), .B(_abc_3927_n504_1), .Y(_abc_3927_n505) );
	INVX1 INVX1_21 ( .A(currentrow_10_), .Y(_abc_3927_n506) );
	AND2X2 AND2X2_13 ( .A(_abc_3927_n506), .B(reg_vf_value_10_), .Y(_abc_3927_n507) );
	NAND2X1 NAND2X1_38 ( .A(_abc_3927_n507), .B(_abc_3927_n440_1), .Y(_abc_3927_n508) );
	NAND2X1 NAND2X1_39 ( .A(_abc_3927_n439_1), .B(_abc_3927_n508), .Y(_abc_3927_n509) );
	NOR2X1 NOR2X1_27 ( .A(_abc_3927_n509), .B(_abc_3927_n505), .Y(_abc_3927_n510_1) );
	NOR2X1 NOR2X1_28 ( .A(_abc_3927_n437_1), .B(_abc_3927_n510_1), .Y(_abc_3927_n511) );
	AND2X2 AND2X2_14 ( .A(_abc_3927_n435_1), .B(_abc_3927_n430_1), .Y(_abc_3927_n512) );
	NOR2X1 NOR2X1_29 ( .A(_abc_3927_n434_1), .B(_abc_3927_n512), .Y(_abc_3927_n513_1) );
	NOR2X1 NOR2X1_30 ( .A(_abc_3927_n427_1), .B(_abc_3927_n513_1), .Y(_abc_3927_n514) );
	NAND2X1 NAND2X1_40 ( .A(_abc_3927_n424), .B(_abc_3927_n421), .Y(_abc_3927_n515) );
	NAND2X1 NAND2X1_41 ( .A(_abc_3927_n420), .B(_abc_3927_n515), .Y(_abc_3927_n516_1) );
	OR2X2 OR2X2_12 ( .A(_abc_3927_n514), .B(_abc_3927_n516_1), .Y(_abc_3927_n517) );
	NOR2X1 NOR2X1_31 ( .A(_abc_3927_n511), .B(_abc_3927_n517), .Y(_abc_3927_n518) );
	NAND2X1 NAND2X1_42 ( .A(_abc_3927_n518), .B(_abc_3927_n502), .Y(_abc_3927_n519_1) );
	INVX2 INVX2_14 ( .A(currentcol_15_), .Y(_abc_3927_n520) );
	NAND2X1 NAND2X1_43 ( .A(reg_hf_value_15_), .B(_abc_3927_n520), .Y(_abc_3927_n521_1) );
	OR2X2 OR2X2_13 ( .A(_abc_3927_n520), .B(reg_hf_value_15_), .Y(_abc_3927_n522_1) );
	AND2X2 AND2X2_15 ( .A(_abc_3927_n522_1), .B(_abc_3927_n521_1), .Y(_abc_3927_n523) );
	INVX4 INVX4_1 ( .A(currentcol_14_), .Y(_abc_3927_n524) );
	NOR2X1 NOR2X1_32 ( .A(reg_hf_value_14_), .B(_abc_3927_n524), .Y(_abc_3927_n525) );
	AND2X2 AND2X2_16 ( .A(_abc_3927_n524), .B(reg_hf_value_14_), .Y(_abc_3927_n526) );
	NOR2X1 NOR2X1_33 ( .A(_abc_3927_n525), .B(_abc_3927_n526), .Y(_abc_3927_n527_1) );
	NAND2X1 NAND2X1_44 ( .A(_abc_3927_n527_1), .B(_abc_3927_n523), .Y(_abc_3927_n528) );
	INVX2 INVX2_15 ( .A(currentcol_13_), .Y(_abc_3927_n529) );
	NAND2X1 NAND2X1_45 ( .A(reg_hf_value_13_), .B(_abc_3927_n529), .Y(_abc_3927_n530) );
	INVX2 INVX2_16 ( .A(currentcol_12_), .Y(_abc_3927_n531) );
	NAND2X1 NAND2X1_46 ( .A(reg_hf_value_12_), .B(_abc_3927_n531), .Y(_abc_3927_n532) );
	NAND2X1 NAND2X1_47 ( .A(_abc_3927_n530), .B(_abc_3927_n532), .Y(_abc_3927_n533) );
	OR2X2 OR2X2_14 ( .A(_abc_3927_n529), .B(reg_hf_value_13_), .Y(_abc_3927_n534) );
	OR2X2 OR2X2_15 ( .A(_abc_3927_n531), .B(reg_hf_value_12_), .Y(_abc_3927_n535) );
	NAND2X1 NAND2X1_48 ( .A(_abc_3927_n534), .B(_abc_3927_n535), .Y(_abc_3927_n536) );
	OR2X2 OR2X2_16 ( .A(_abc_3927_n536), .B(_abc_3927_n533), .Y(_abc_3927_n537) );
	NOR2X1 NOR2X1_34 ( .A(_abc_3927_n528), .B(_abc_3927_n537), .Y(_abc_3927_n538) );
	INVX2 INVX2_17 ( .A(currentcol_11_), .Y(_abc_3927_n539) );
	NAND2X1 NAND2X1_49 ( .A(reg_hf_value_11_), .B(_abc_3927_n539), .Y(_abc_3927_n540) );
	INVX1 INVX1_22 ( .A(reg_hf_value_11_), .Y(_abc_3927_n541) );
	NAND2X1 NAND2X1_50 ( .A(currentcol_11_), .B(_abc_3927_n541), .Y(_abc_3927_n542) );
	AND2X2 AND2X2_17 ( .A(_abc_3927_n540), .B(_abc_3927_n542), .Y(_abc_3927_n543) );
	XNOR2X1 XNOR2X1_11 ( .A(currentcol_10_), .B(reg_hf_value_10_), .Y(_abc_3927_n544) );
	NAND2X1 NAND2X1_51 ( .A(_abc_3927_n544), .B(_abc_3927_n543), .Y(_abc_3927_n545) );
	INVX2 INVX2_18 ( .A(currentcol_9_), .Y(_abc_3927_n546) );
	NAND2X1 NAND2X1_52 ( .A(reg_hf_value_9_), .B(_abc_3927_n546), .Y(_abc_3927_n547) );
	INVX2 INVX2_19 ( .A(currentcol_8_), .Y(_abc_3927_n548) );
	NAND2X1 NAND2X1_53 ( .A(reg_hf_value_8_), .B(_abc_3927_n548), .Y(_abc_3927_n549) );
	NAND2X1 NAND2X1_54 ( .A(_abc_3927_n547), .B(_abc_3927_n549), .Y(_abc_3927_n550) );
	NOR2X1 NOR2X1_35 ( .A(reg_hf_value_8_), .B(_abc_3927_n548), .Y(_abc_3927_n551) );
	NOR2X1 NOR2X1_36 ( .A(reg_hf_value_9_), .B(_abc_3927_n546), .Y(_abc_3927_n552) );
	OR2X2 OR2X2_17 ( .A(_abc_3927_n551), .B(_abc_3927_n552), .Y(_abc_3927_n553) );
	OR2X2 OR2X2_18 ( .A(_abc_3927_n553), .B(_abc_3927_n550), .Y(_abc_3927_n554) );
	NOR2X1 NOR2X1_37 ( .A(_abc_3927_n545), .B(_abc_3927_n554), .Y(_abc_3927_n555) );
	AND2X2 AND2X2_18 ( .A(_abc_3927_n555), .B(_abc_3927_n538), .Y(_abc_3927_n556) );
	INVX1 INVX1_23 ( .A(reg_hf_value_7_), .Y(_abc_3927_n557) );
	NAND2X1 NAND2X1_55 ( .A(currentcol_7_), .B(_abc_3927_n557), .Y(_abc_3927_n558) );
	NOR2X1 NOR2X1_38 ( .A(currentcol_7_), .B(_abc_3927_n557), .Y(_abc_3927_n559) );
	INVX1 INVX1_24 ( .A(_abc_3927_n559), .Y(_abc_3927_n560) );
	AND2X2 AND2X2_19 ( .A(_abc_3927_n560), .B(_abc_3927_n558), .Y(_abc_3927_n561) );
	INVX2 INVX2_20 ( .A(currentcol_6_), .Y(_abc_3927_n562) );
	NOR2X1 NOR2X1_39 ( .A(reg_hf_value_6_), .B(_abc_3927_n562), .Y(_abc_3927_n563) );
	AND2X2 AND2X2_20 ( .A(_abc_3927_n562), .B(reg_hf_value_6_), .Y(_abc_3927_n564) );
	NOR2X1 NOR2X1_40 ( .A(_abc_3927_n563), .B(_abc_3927_n564), .Y(_abc_3927_n565) );
	NAND2X1 NAND2X1_56 ( .A(_abc_3927_n565), .B(_abc_3927_n561), .Y(_abc_3927_n566) );
	INVX2 INVX2_21 ( .A(currentcol_5_), .Y(_abc_3927_n567) );
	NAND2X1 NAND2X1_57 ( .A(reg_hf_value_5_), .B(_abc_3927_n567), .Y(_abc_3927_n568) );
	INVX2 INVX2_22 ( .A(currentcol_4_), .Y(_abc_3927_n569) );
	NAND2X1 NAND2X1_58 ( .A(reg_hf_value_4_), .B(_abc_3927_n569), .Y(_abc_3927_n570) );
	NAND2X1 NAND2X1_59 ( .A(_abc_3927_n568), .B(_abc_3927_n570), .Y(_abc_3927_n571) );
	OR2X2 OR2X2_19 ( .A(_abc_3927_n567), .B(reg_hf_value_5_), .Y(_abc_3927_n572) );
	OR2X2 OR2X2_20 ( .A(_abc_3927_n569), .B(reg_hf_value_4_), .Y(_abc_3927_n573) );
	NAND2X1 NAND2X1_60 ( .A(_abc_3927_n572), .B(_abc_3927_n573), .Y(_abc_3927_n574) );
	OR2X2 OR2X2_21 ( .A(_abc_3927_n574), .B(_abc_3927_n571), .Y(_abc_3927_n575) );
	NOR2X1 NOR2X1_41 ( .A(_abc_3927_n575), .B(_abc_3927_n566), .Y(_abc_3927_n576) );
	INVX2 INVX2_23 ( .A(currentcol_3_), .Y(_abc_3927_n577) );
	NAND2X1 NAND2X1_61 ( .A(reg_hf_value_3_), .B(_abc_3927_n577), .Y(_abc_3927_n578) );
	OR2X2 OR2X2_22 ( .A(_abc_3927_n577), .B(reg_hf_value_3_), .Y(_abc_3927_n579) );
	NAND2X1 NAND2X1_62 ( .A(_abc_3927_n578), .B(_abc_3927_n579), .Y(_abc_3927_n580) );
	XOR2X1 XOR2X1_11 ( .A(currentcol_2_), .B(reg_hf_value_2_), .Y(_abc_3927_n581) );
	NOR2X1 NOR2X1_42 ( .A(_abc_3927_n581), .B(_abc_3927_n580), .Y(_abc_3927_n582) );
	INVX2 INVX2_24 ( .A(currentcol_1_), .Y(_abc_3927_n583) );
	NAND2X1 NAND2X1_63 ( .A(reg_hf_value_1_), .B(_abc_3927_n583), .Y(_abc_3927_n584) );
	INVX2 INVX2_25 ( .A(currentcol_0_), .Y(_abc_3927_n585) );
	OR2X2 OR2X2_23 ( .A(_abc_3927_n585), .B(reg_hf_value_0_), .Y(_abc_3927_n586) );
	XNOR2X1 XNOR2X1_12 ( .A(currentcol_1_), .B(reg_hf_value_1_), .Y(_abc_3927_n587) );
	NAND2X1 NAND2X1_64 ( .A(_abc_3927_n586), .B(_abc_3927_n587), .Y(_abc_3927_n588) );
	NAND2X1 NAND2X1_65 ( .A(_abc_3927_n584), .B(_abc_3927_n588), .Y(_abc_3927_n589) );
	NAND2X1 NAND2X1_66 ( .A(_abc_3927_n582), .B(_abc_3927_n589), .Y(_abc_3927_n590) );
	INVX1 INVX1_25 ( .A(currentcol_2_), .Y(_abc_3927_n591) );
	AND2X2 AND2X2_21 ( .A(_abc_3927_n591), .B(reg_hf_value_2_), .Y(_abc_3927_n592) );
	NAND2X1 NAND2X1_67 ( .A(_abc_3927_n592), .B(_abc_3927_n579), .Y(_abc_3927_n593) );
	AND2X2 AND2X2_22 ( .A(_abc_3927_n593), .B(_abc_3927_n578), .Y(_abc_3927_n594) );
	NAND2X1 NAND2X1_68 ( .A(_abc_3927_n594), .B(_abc_3927_n590), .Y(_abc_3927_n595) );
	NAND2X1 NAND2X1_69 ( .A(_abc_3927_n576), .B(_abc_3927_n595), .Y(_abc_3927_n596) );
	NAND2X1 NAND2X1_70 ( .A(_abc_3927_n558), .B(_abc_3927_n564), .Y(_abc_3927_n597) );
	NAND2X1 NAND2X1_71 ( .A(_abc_3927_n560), .B(_abc_3927_n597), .Y(_abc_3927_n598) );
	NAND2X1 NAND2X1_72 ( .A(_abc_3927_n572), .B(_abc_3927_n571), .Y(_abc_3927_n599) );
	NOR2X1 NOR2X1_43 ( .A(_abc_3927_n599), .B(_abc_3927_n566), .Y(_abc_3927_n600) );
	NOR2X1 NOR2X1_44 ( .A(_abc_3927_n598), .B(_abc_3927_n600), .Y(_abc_3927_n601) );
	NAND2X1 NAND2X1_73 ( .A(_abc_3927_n596), .B(_abc_3927_n601), .Y(_abc_3927_n602) );
	NAND2X1 NAND2X1_74 ( .A(_abc_3927_n556), .B(_abc_3927_n602), .Y(_abc_3927_n603) );
	INVX2 INVX2_26 ( .A(currentcol_10_), .Y(_abc_3927_n604) );
	NAND2X1 NAND2X1_75 ( .A(reg_hf_value_10_), .B(_abc_3927_n604), .Y(_abc_3927_n605) );
	NAND2X1 NAND2X1_76 ( .A(_abc_3927_n540), .B(_abc_3927_n605), .Y(_abc_3927_n606) );
	NAND2X1 NAND2X1_77 ( .A(_abc_3927_n542), .B(_abc_3927_n606), .Y(_abc_3927_n607) );
	NOR2X1 NOR2X1_45 ( .A(_abc_3927_n552), .B(_abc_3927_n545), .Y(_abc_3927_n608) );
	NAND2X1 NAND2X1_78 ( .A(_abc_3927_n550), .B(_abc_3927_n608), .Y(_abc_3927_n609) );
	NAND2X1 NAND2X1_79 ( .A(_abc_3927_n607), .B(_abc_3927_n609), .Y(_abc_3927_n610) );
	NAND2X1 NAND2X1_80 ( .A(_abc_3927_n538), .B(_abc_3927_n610), .Y(_abc_3927_n611) );
	NAND2X1 NAND2X1_81 ( .A(_abc_3927_n526), .B(_abc_3927_n522_1), .Y(_abc_3927_n612) );
	NAND2X1 NAND2X1_82 ( .A(_abc_3927_n521_1), .B(_abc_3927_n612), .Y(_abc_3927_n613) );
	NAND2X1 NAND2X1_83 ( .A(_abc_3927_n534), .B(_abc_3927_n533), .Y(_abc_3927_n614_1) );
	NOR2X1 NOR2X1_46 ( .A(_abc_3927_n614_1), .B(_abc_3927_n528), .Y(_abc_3927_n615) );
	NOR2X1 NOR2X1_47 ( .A(_abc_3927_n613), .B(_abc_3927_n615), .Y(_abc_3927_n616) );
	AND2X2 AND2X2_23 ( .A(_abc_3927_n611), .B(_abc_3927_n616), .Y(_abc_3927_n617) );
	NAND2X1 NAND2X1_84 ( .A(_abc_3927_n603), .B(_abc_3927_n617), .Y(_abc_3927_n618) );
	NAND2X1 NAND2X1_85 ( .A(reg_hf_value_0_), .B(_abc_3927_n585), .Y(_abc_3927_n619_1) );
	NAND2X1 NAND2X1_86 ( .A(_abc_3927_n619_1), .B(_abc_3927_n582), .Y(_abc_3927_n620) );
	NOR2X1 NOR2X1_48 ( .A(_abc_3927_n588), .B(_abc_3927_n620), .Y(_abc_3927_n621_1) );
	AND2X2 AND2X2_24 ( .A(_abc_3927_n621_1), .B(_abc_3927_n576), .Y(_abc_3927_n622_1) );
	AND2X2 AND2X2_25 ( .A(_abc_3927_n622_1), .B(_abc_3927_n556), .Y(_abc_3927_n623) );
	NAND2X1 NAND2X1_87 ( .A(reg_vf_value_0_), .B(_abc_3927_n480_1), .Y(_abc_3927_n624) );
	NAND2X1 NAND2X1_88 ( .A(_abc_3927_n624), .B(_abc_3927_n477), .Y(_abc_3927_n625) );
	NOR2X1 NOR2X1_49 ( .A(_abc_3927_n483_1), .B(_abc_3927_n625), .Y(_abc_3927_n626_1) );
	NAND2X1 NAND2X1_89 ( .A(_abc_3927_n471), .B(_abc_3927_n626_1), .Y(_abc_3927_n627_1) );
	NOR2X1 NOR2X1_50 ( .A(_abc_3927_n627_1), .B(_abc_3927_n455), .Y(_abc_3927_n628) );
	NOR2X1 NOR2X1_51 ( .A(_abc_3927_n628), .B(_abc_3927_n623), .Y(_abc_3927_n629) );
	AND2X2 AND2X2_26 ( .A(_abc_3927_n629), .B(_abc_3927_n618), .Y(_abc_3927_n630_1) );
	NAND2X1 NAND2X1_90 ( .A(_abc_3927_n519_1), .B(_abc_3927_n630_1), .Y(_abc_3927_n631) );
	NAND2X1 NAND2X1_91 ( .A(reg_hv_value_15_), .B(_abc_3927_n520), .Y(_abc_3927_n632_1) );
	OR2X2 OR2X2_24 ( .A(_abc_3927_n520), .B(reg_hv_value_15_), .Y(_abc_3927_n633) );
	AND2X2 AND2X2_27 ( .A(_abc_3927_n633), .B(_abc_3927_n632_1), .Y(_abc_3927_n634_1) );
	NOR2X1 NOR2X1_52 ( .A(reg_hv_value_14_), .B(_abc_3927_n524), .Y(_abc_3927_n635) );
	AND2X2 AND2X2_28 ( .A(_abc_3927_n524), .B(reg_hv_value_14_), .Y(_abc_3927_n636_1) );
	NOR2X1 NOR2X1_53 ( .A(_abc_3927_n635), .B(_abc_3927_n636_1), .Y(_abc_3927_n637) );
	NAND2X1 NAND2X1_92 ( .A(_abc_3927_n637), .B(_abc_3927_n634_1), .Y(_abc_3927_n638_1) );
	NAND2X1 NAND2X1_93 ( .A(reg_hv_value_13_), .B(_abc_3927_n529), .Y(_abc_3927_n639) );
	NAND2X1 NAND2X1_94 ( .A(reg_hv_value_12_), .B(_abc_3927_n531), .Y(_abc_3927_n640_1) );
	NAND2X1 NAND2X1_95 ( .A(_abc_3927_n639), .B(_abc_3927_n640_1), .Y(_abc_3927_n641) );
	OR2X2 OR2X2_25 ( .A(_abc_3927_n529), .B(reg_hv_value_13_), .Y(_abc_3927_n642_1) );
	OR2X2 OR2X2_26 ( .A(_abc_3927_n531), .B(reg_hv_value_12_), .Y(_abc_3927_n643) );
	NAND2X1 NAND2X1_96 ( .A(_abc_3927_n642_1), .B(_abc_3927_n643), .Y(_abc_3927_n644_1) );
	OR2X2 OR2X2_27 ( .A(_abc_3927_n644_1), .B(_abc_3927_n641), .Y(_abc_3927_n645) );
	NOR2X1 NOR2X1_54 ( .A(_abc_3927_n638_1), .B(_abc_3927_n645), .Y(_abc_3927_n646_1) );
	NAND2X1 NAND2X1_97 ( .A(reg_hv_value_11_), .B(_abc_3927_n539), .Y(_abc_3927_n647) );
	NAND2X1 NAND2X1_98 ( .A(reg_hv_value_10_), .B(_abc_3927_n604), .Y(_abc_3927_n648_1) );
	NAND2X1 NAND2X1_99 ( .A(_abc_3927_n647), .B(_abc_3927_n648_1), .Y(_abc_3927_n649) );
	OR2X2 OR2X2_28 ( .A(_abc_3927_n539), .B(reg_hv_value_11_), .Y(_abc_3927_n650_1) );
	OR2X2 OR2X2_29 ( .A(_abc_3927_n604), .B(reg_hv_value_10_), .Y(_abc_3927_n651) );
	NAND2X1 NAND2X1_100 ( .A(_abc_3927_n650_1), .B(_abc_3927_n651), .Y(_abc_3927_n652_1) );
	NOR2X1 NOR2X1_55 ( .A(_abc_3927_n649), .B(_abc_3927_n652_1), .Y(_abc_3927_n653) );
	NAND2X1 NAND2X1_101 ( .A(reg_hv_value_9_), .B(_abc_3927_n546), .Y(_abc_3927_n654_1) );
	NAND2X1 NAND2X1_102 ( .A(reg_hv_value_8_), .B(_abc_3927_n548), .Y(_abc_3927_n655) );
	NAND2X1 NAND2X1_103 ( .A(_abc_3927_n654_1), .B(_abc_3927_n655), .Y(_abc_3927_n656_1) );
	OR2X2 OR2X2_30 ( .A(_abc_3927_n548), .B(reg_hv_value_8_), .Y(_abc_3927_n657) );
	OR2X2 OR2X2_31 ( .A(_abc_3927_n546), .B(reg_hv_value_9_), .Y(_abc_3927_n658_1) );
	NAND2X1 NAND2X1_104 ( .A(_abc_3927_n657), .B(_abc_3927_n658_1), .Y(_abc_3927_n659) );
	NOR2X1 NOR2X1_56 ( .A(_abc_3927_n656_1), .B(_abc_3927_n659), .Y(_abc_3927_n660) );
	AND2X2 AND2X2_29 ( .A(_abc_3927_n653), .B(_abc_3927_n660), .Y(_abc_3927_n661) );
	AND2X2 AND2X2_30 ( .A(_abc_3927_n646_1), .B(_abc_3927_n661), .Y(_abc_3927_n662) );
	INVX2 INVX2_27 ( .A(currentcol_7_), .Y(_abc_3927_n663) );
	NAND2X1 NAND2X1_105 ( .A(reg_hv_value_7_), .B(_abc_3927_n663), .Y(_abc_3927_n664) );
	NAND2X1 NAND2X1_106 ( .A(reg_hv_value_6_), .B(_abc_3927_n562), .Y(_abc_3927_n665) );
	NAND2X1 NAND2X1_107 ( .A(_abc_3927_n664), .B(_abc_3927_n665), .Y(_abc_3927_n666) );
	NOR2X1 NOR2X1_57 ( .A(reg_hv_value_7_), .B(_abc_3927_n663), .Y(_abc_3927_n667) );
	NOR2X1 NOR2X1_58 ( .A(reg_hv_value_6_), .B(_abc_3927_n562), .Y(_abc_3927_n668) );
	OR2X2 OR2X2_32 ( .A(_abc_3927_n667), .B(_abc_3927_n668), .Y(_abc_3927_n669) );
	OR2X2 OR2X2_33 ( .A(_abc_3927_n669), .B(_abc_3927_n666), .Y(_abc_3927_n670) );
	NAND2X1 NAND2X1_108 ( .A(reg_hv_value_5_), .B(_abc_3927_n567), .Y(_abc_3927_n671_1) );
	NAND2X1 NAND2X1_109 ( .A(reg_hv_value_4_), .B(_abc_3927_n569), .Y(_abc_3927_n672) );
	NAND2X1 NAND2X1_110 ( .A(_abc_3927_n671_1), .B(_abc_3927_n672), .Y(_abc_3927_n673) );
	OR2X2 OR2X2_34 ( .A(_abc_3927_n567), .B(reg_hv_value_5_), .Y(_abc_3927_n674_1) );
	OR2X2 OR2X2_35 ( .A(_abc_3927_n569), .B(reg_hv_value_4_), .Y(_abc_3927_n675) );
	AND2X2 AND2X2_31 ( .A(_abc_3927_n674_1), .B(_abc_3927_n675), .Y(_abc_3927_n676) );
	INVX1 INVX1_26 ( .A(_abc_3927_n676), .Y(_abc_3927_n677) );
	OR2X2 OR2X2_36 ( .A(_abc_3927_n677), .B(_abc_3927_n673), .Y(_abc_3927_n678) );
	NOR2X1 NOR2X1_59 ( .A(_abc_3927_n670), .B(_abc_3927_n678), .Y(_abc_3927_n679) );
	NAND2X1 NAND2X1_111 ( .A(reg_hv_value_3_), .B(_abc_3927_n577), .Y(_abc_3927_n680) );
	OR2X2 OR2X2_37 ( .A(_abc_3927_n577), .B(reg_hv_value_3_), .Y(_abc_3927_n681) );
	NAND2X1 NAND2X1_112 ( .A(_abc_3927_n680), .B(_abc_3927_n681), .Y(_abc_3927_n682_1) );
	XOR2X1 XOR2X1_12 ( .A(currentcol_2_), .B(reg_hv_value_2_), .Y(_abc_3927_n683_1) );
	NOR2X1 NOR2X1_60 ( .A(_abc_3927_n683_1), .B(_abc_3927_n682_1), .Y(_abc_3927_n684) );
	NAND2X1 NAND2X1_113 ( .A(reg_hv_value_1_), .B(_abc_3927_n583), .Y(_abc_3927_n685_1) );
	INVX1 INVX1_27 ( .A(reg_hv_value_0_), .Y(_abc_3927_n686) );
	NAND2X1 NAND2X1_114 ( .A(currentcol_0_), .B(_abc_3927_n686), .Y(_abc_3927_n687_1) );
	XNOR2X1 XNOR2X1_13 ( .A(currentcol_1_), .B(reg_hv_value_1_), .Y(_abc_3927_n688_1) );
	NAND2X1 NAND2X1_115 ( .A(_abc_3927_n687_1), .B(_abc_3927_n688_1), .Y(_abc_3927_n689_1) );
	NAND2X1 NAND2X1_116 ( .A(_abc_3927_n685_1), .B(_abc_3927_n689_1), .Y(_abc_3927_n690) );
	NAND2X1 NAND2X1_117 ( .A(_abc_3927_n684), .B(_abc_3927_n690), .Y(_abc_3927_n691) );
	AND2X2 AND2X2_32 ( .A(_abc_3927_n591), .B(reg_hv_value_2_), .Y(_abc_3927_n692) );
	NAND2X1 NAND2X1_118 ( .A(_abc_3927_n692), .B(_abc_3927_n681), .Y(_abc_3927_n693) );
	AND2X2 AND2X2_33 ( .A(_abc_3927_n693), .B(_abc_3927_n680), .Y(_abc_3927_n694) );
	NAND2X1 NAND2X1_119 ( .A(_abc_3927_n694), .B(_abc_3927_n691), .Y(_abc_3927_n695) );
	NAND2X1 NAND2X1_120 ( .A(_abc_3927_n695), .B(_abc_3927_n679), .Y(_abc_3927_n696) );
	INVX1 INVX1_28 ( .A(_abc_3927_n667), .Y(_abc_3927_n697) );
	AND2X2 AND2X2_34 ( .A(_abc_3927_n697), .B(_abc_3927_n666), .Y(_abc_3927_n698) );
	NAND2X1 NAND2X1_121 ( .A(_abc_3927_n674_1), .B(_abc_3927_n673), .Y(_abc_3927_n699) );
	NOR2X1 NOR2X1_61 ( .A(_abc_3927_n699), .B(_abc_3927_n670), .Y(_abc_3927_n700) );
	NOR2X1 NOR2X1_62 ( .A(_abc_3927_n698), .B(_abc_3927_n700), .Y(_abc_3927_n701) );
	NAND2X1 NAND2X1_122 ( .A(_abc_3927_n701), .B(_abc_3927_n696), .Y(_abc_3927_n702) );
	NAND2X1 NAND2X1_123 ( .A(_abc_3927_n662), .B(_abc_3927_n702), .Y(_abc_3927_n703) );
	NAND2X1 NAND2X1_124 ( .A(_abc_3927_n650_1), .B(_abc_3927_n649), .Y(_abc_3927_n704) );
	AND2X2 AND2X2_35 ( .A(_abc_3927_n656_1), .B(_abc_3927_n658_1), .Y(_abc_3927_n705) );
	NAND2X1 NAND2X1_125 ( .A(_abc_3927_n705), .B(_abc_3927_n653), .Y(_abc_3927_n706) );
	NAND2X1 NAND2X1_126 ( .A(_abc_3927_n704), .B(_abc_3927_n706), .Y(_abc_3927_n707) );
	NAND2X1 NAND2X1_127 ( .A(_abc_3927_n646_1), .B(_abc_3927_n707), .Y(_abc_3927_n708) );
	NAND2X1 NAND2X1_128 ( .A(_abc_3927_n636_1), .B(_abc_3927_n633), .Y(_abc_3927_n709) );
	NAND2X1 NAND2X1_129 ( .A(_abc_3927_n632_1), .B(_abc_3927_n709), .Y(_abc_3927_n710) );
	NAND2X1 NAND2X1_130 ( .A(_abc_3927_n642_1), .B(_abc_3927_n641), .Y(_abc_3927_n711) );
	NOR2X1 NOR2X1_63 ( .A(_abc_3927_n711), .B(_abc_3927_n638_1), .Y(_abc_3927_n712) );
	NOR2X1 NOR2X1_64 ( .A(_abc_3927_n710), .B(_abc_3927_n712), .Y(_abc_3927_n713) );
	AND2X2 AND2X2_36 ( .A(_abc_3927_n708), .B(_abc_3927_n713), .Y(_abc_3927_n714) );
	NAND2X1 NAND2X1_131 ( .A(_abc_3927_n714), .B(_abc_3927_n703), .Y(_abc_3927_n715) );
	NAND2X1 NAND2X1_132 ( .A(reg_hv_value_0_), .B(_abc_3927_n585), .Y(_abc_3927_n716) );
	NAND2X1 NAND2X1_133 ( .A(_abc_3927_n716), .B(_abc_3927_n684), .Y(_abc_3927_n717) );
	NOR2X1 NOR2X1_65 ( .A(_abc_3927_n689_1), .B(_abc_3927_n717), .Y(_abc_3927_n718) );
	AND2X2 AND2X2_37 ( .A(_abc_3927_n679), .B(_abc_3927_n718), .Y(_abc_3927_n719) );
	NAND2X1 NAND2X1_134 ( .A(_abc_3927_n662), .B(_abc_3927_n719), .Y(_abc_3927_n720) );
	NAND2X1 NAND2X1_135 ( .A(_abc_3927_n720), .B(_abc_3927_n715), .Y(_abc_3927_n721) );
	NAND2X1 NAND2X1_136 ( .A(reg_vv_value_15_), .B(_abc_3927_n419), .Y(_abc_3927_n722) );
	OR2X2 OR2X2_38 ( .A(_abc_3927_n419), .B(reg_vv_value_15_), .Y(_abc_3927_n723) );
	AND2X2 AND2X2_38 ( .A(_abc_3927_n723), .B(_abc_3927_n722), .Y(_abc_3927_n724) );
	AND2X2 AND2X2_39 ( .A(_abc_3927_n423), .B(reg_vv_value_14_), .Y(_abc_3927_n725) );
	NOR2X1 NOR2X1_66 ( .A(reg_vv_value_14_), .B(_abc_3927_n423), .Y(_abc_3927_n726) );
	NOR2X1 NOR2X1_67 ( .A(_abc_3927_n726), .B(_abc_3927_n725), .Y(_abc_3927_n727) );
	NAND2X1 NAND2X1_137 ( .A(_abc_3927_n727), .B(_abc_3927_n724), .Y(_abc_3927_n728) );
	NOR2X1 NOR2X1_68 ( .A(reg_vv_value_12_), .B(_abc_3927_n428_1), .Y(_abc_3927_n729) );
	AND2X2 AND2X2_40 ( .A(_abc_3927_n428_1), .B(reg_vv_value_12_), .Y(_abc_3927_n730) );
	NOR2X1 NOR2X1_69 ( .A(_abc_3927_n729), .B(_abc_3927_n730), .Y(_abc_3927_n731) );
	OR2X2 OR2X2_39 ( .A(_abc_3927_n432_1), .B(reg_vv_value_13_), .Y(_abc_3927_n732) );
	NAND2X1 NAND2X1_138 ( .A(reg_vv_value_13_), .B(_abc_3927_n432_1), .Y(_abc_3927_n733) );
	AND2X2 AND2X2_41 ( .A(_abc_3927_n732), .B(_abc_3927_n733), .Y(_abc_3927_n734) );
	NAND2X1 NAND2X1_139 ( .A(_abc_3927_n731), .B(_abc_3927_n734), .Y(_abc_3927_n735) );
	NOR2X1 NOR2X1_70 ( .A(_abc_3927_n728), .B(_abc_3927_n735), .Y(_abc_3927_n736) );
	NAND2X1 NAND2X1_140 ( .A(reg_vv_value_11_), .B(_abc_3927_n438_1), .Y(_abc_3927_n737) );
	OR2X2 OR2X2_40 ( .A(_abc_3927_n438_1), .B(reg_vv_value_11_), .Y(_abc_3927_n738) );
	NAND2X1 NAND2X1_141 ( .A(_abc_3927_n737), .B(_abc_3927_n738), .Y(_abc_3927_n739) );
	XOR2X1 XOR2X1_13 ( .A(reg_vv_value_10_), .B(currentrow_10_), .Y(_abc_3927_n740) );
	NOR2X1 NOR2X1_71 ( .A(_abc_3927_n740), .B(_abc_3927_n739), .Y(_abc_3927_n741) );
	INVX1 INVX1_29 ( .A(currentrow_8_), .Y(_abc_3927_n742) );
	NAND2X1 NAND2X1_142 ( .A(reg_vv_value_8_), .B(_abc_3927_n742), .Y(_abc_3927_n743) );
	NAND2X1 NAND2X1_143 ( .A(reg_vv_value_9_), .B(_abc_3927_n446), .Y(_abc_3927_n744) );
	NAND2X1 NAND2X1_144 ( .A(_abc_3927_n743), .B(_abc_3927_n744), .Y(_abc_3927_n745) );
	OR2X2 OR2X2_41 ( .A(_abc_3927_n742), .B(reg_vv_value_8_), .Y(_abc_3927_n746) );
	OR2X2 OR2X2_42 ( .A(_abc_3927_n446), .B(reg_vv_value_9_), .Y(_abc_3927_n747) );
	NAND2X1 NAND2X1_145 ( .A(_abc_3927_n746), .B(_abc_3927_n747), .Y(_abc_3927_n748) );
	NOR2X1 NOR2X1_72 ( .A(_abc_3927_n745), .B(_abc_3927_n748), .Y(_abc_3927_n749) );
	AND2X2 AND2X2_42 ( .A(_abc_3927_n749), .B(_abc_3927_n741), .Y(_abc_3927_n750) );
	AND2X2 AND2X2_43 ( .A(_abc_3927_n736), .B(_abc_3927_n750), .Y(_abc_3927_n751) );
	NAND2X1 NAND2X1_146 ( .A(reg_vv_value_7_), .B(_abc_3927_n456), .Y(_abc_3927_n752) );
	OR2X2 OR2X2_43 ( .A(_abc_3927_n456), .B(reg_vv_value_7_), .Y(_abc_3927_n753) );
	NAND2X1 NAND2X1_147 ( .A(_abc_3927_n752), .B(_abc_3927_n753), .Y(_abc_3927_n754) );
	XOR2X1 XOR2X1_14 ( .A(reg_vv_value_6_), .B(currentrow_6_), .Y(_abc_3927_n755) );
	NOR2X1 NOR2X1_73 ( .A(_abc_3927_n755), .B(_abc_3927_n754), .Y(_abc_3927_n756) );
	INVX1 INVX1_30 ( .A(_abc_3927_n756), .Y(_abc_3927_n757) );
	XNOR2X1 XNOR2X1_14 ( .A(reg_vv_value_5_), .B(currentrow_5_), .Y(_abc_3927_n758) );
	XNOR2X1 XNOR2X1_15 ( .A(reg_vv_value_4_), .B(currentrow_4_), .Y(_abc_3927_n759) );
	NAND2X1 NAND2X1_148 ( .A(_abc_3927_n758), .B(_abc_3927_n759), .Y(_abc_3927_n760) );
	NOR2X1 NOR2X1_74 ( .A(_abc_3927_n760), .B(_abc_3927_n757), .Y(_abc_3927_n761) );
	NAND2X1 NAND2X1_149 ( .A(reg_vv_value_3_), .B(_abc_3927_n472), .Y(_abc_3927_n762) );
	OR2X2 OR2X2_44 ( .A(_abc_3927_n472), .B(reg_vv_value_3_), .Y(_abc_3927_n763) );
	NAND2X1 NAND2X1_150 ( .A(_abc_3927_n762), .B(_abc_3927_n763), .Y(_abc_3927_n764) );
	XOR2X1 XOR2X1_15 ( .A(reg_vv_value_2_), .B(currentrow_2_), .Y(_abc_3927_n765) );
	NOR2X1 NOR2X1_75 ( .A(_abc_3927_n765), .B(_abc_3927_n764), .Y(_abc_3927_n766) );
	AND2X2 AND2X2_44 ( .A(_abc_3927_n478_1), .B(reg_vv_value_1_), .Y(_abc_3927_n767) );
	INVX1 INVX1_31 ( .A(_abc_3927_n767), .Y(_abc_3927_n768) );
	OR2X2 OR2X2_45 ( .A(_abc_3927_n480_1), .B(reg_vv_value_0_), .Y(_abc_3927_n769) );
	NOR2X1 NOR2X1_76 ( .A(reg_vv_value_1_), .B(_abc_3927_n478_1), .Y(_abc_3927_n770) );
	NOR2X1 NOR2X1_77 ( .A(_abc_3927_n770), .B(_abc_3927_n767), .Y(_abc_3927_n771) );
	NAND2X1 NAND2X1_151 ( .A(_abc_3927_n769), .B(_abc_3927_n771), .Y(_abc_3927_n772) );
	NAND2X1 NAND2X1_152 ( .A(_abc_3927_n768), .B(_abc_3927_n772), .Y(_abc_3927_n773) );
	NAND2X1 NAND2X1_153 ( .A(_abc_3927_n766), .B(_abc_3927_n773), .Y(_abc_3927_n774) );
	AND2X2 AND2X2_45 ( .A(_abc_3927_n486_1), .B(reg_vv_value_2_), .Y(_abc_3927_n775) );
	NAND2X1 NAND2X1_154 ( .A(_abc_3927_n775), .B(_abc_3927_n763), .Y(_abc_3927_n776) );
	AND2X2 AND2X2_46 ( .A(_abc_3927_n776), .B(_abc_3927_n762), .Y(_abc_3927_n777) );
	NAND2X1 NAND2X1_155 ( .A(_abc_3927_n777), .B(_abc_3927_n774), .Y(_abc_3927_n778) );
	NAND2X1 NAND2X1_156 ( .A(_abc_3927_n761), .B(_abc_3927_n778), .Y(_abc_3927_n779_1) );
	NAND2X1 NAND2X1_157 ( .A(reg_vv_value_5_), .B(_abc_3927_n462), .Y(_abc_3927_n780_1) );
	AND2X2 AND2X2_47 ( .A(_abc_3927_n464), .B(reg_vv_value_4_), .Y(_abc_3927_n781_1) );
	NAND2X1 NAND2X1_158 ( .A(_abc_3927_n781_1), .B(_abc_3927_n758), .Y(_abc_3927_n782_1) );
	NAND2X1 NAND2X1_159 ( .A(_abc_3927_n780_1), .B(_abc_3927_n782_1), .Y(_abc_3927_n783_1) );
	AND2X2 AND2X2_48 ( .A(_abc_3927_n783_1), .B(_abc_3927_n756), .Y(_abc_3927_n784_1) );
	AND2X2 AND2X2_49 ( .A(_abc_3927_n496), .B(reg_vv_value_6_), .Y(_abc_3927_n785_1) );
	NAND2X1 NAND2X1_160 ( .A(_abc_3927_n785_1), .B(_abc_3927_n753), .Y(_abc_3927_n786_1) );
	NAND2X1 NAND2X1_161 ( .A(_abc_3927_n752), .B(_abc_3927_n786_1), .Y(_abc_3927_n787_1) );
	NOR2X1 NOR2X1_78 ( .A(_abc_3927_n787_1), .B(_abc_3927_n784_1), .Y(_abc_3927_n788_1) );
	NAND2X1 NAND2X1_162 ( .A(_abc_3927_n788_1), .B(_abc_3927_n779_1), .Y(_abc_3927_n789_1) );
	NAND2X1 NAND2X1_163 ( .A(_abc_3927_n751), .B(_abc_3927_n789_1), .Y(_abc_3927_n790_1) );
	INVX1 INVX1_32 ( .A(_abc_3927_n743), .Y(_abc_3927_n791_1) );
	NAND2X1 NAND2X1_164 ( .A(_abc_3927_n747), .B(_abc_3927_n791_1), .Y(_abc_3927_n792_1) );
	NAND2X1 NAND2X1_165 ( .A(_abc_3927_n744), .B(_abc_3927_n792_1), .Y(_abc_3927_n793_1) );
	NAND2X1 NAND2X1_166 ( .A(_abc_3927_n793_1), .B(_abc_3927_n741), .Y(_abc_3927_n794_1) );
	AND2X2 AND2X2_50 ( .A(_abc_3927_n506), .B(reg_vv_value_10_), .Y(_abc_3927_n795) );
	NAND2X1 NAND2X1_167 ( .A(_abc_3927_n795), .B(_abc_3927_n738), .Y(_abc_3927_n796) );
	AND2X2 AND2X2_51 ( .A(_abc_3927_n796), .B(_abc_3927_n737), .Y(_abc_3927_n797) );
	NAND2X1 NAND2X1_168 ( .A(_abc_3927_n797), .B(_abc_3927_n794_1), .Y(_abc_3927_n798) );
	NAND2X1 NAND2X1_169 ( .A(_abc_3927_n736), .B(_abc_3927_n798), .Y(_abc_3927_n799) );
	NAND2X1 NAND2X1_170 ( .A(_abc_3927_n730), .B(_abc_3927_n732), .Y(_abc_3927_n800) );
	AND2X2 AND2X2_52 ( .A(_abc_3927_n800), .B(_abc_3927_n733), .Y(_abc_3927_n801) );
	NOR2X1 NOR2X1_79 ( .A(_abc_3927_n801), .B(_abc_3927_n728), .Y(_abc_3927_n802) );
	NAND2X1 NAND2X1_171 ( .A(_abc_3927_n725), .B(_abc_3927_n723), .Y(_abc_3927_n803) );
	NAND2X1 NAND2X1_172 ( .A(_abc_3927_n722), .B(_abc_3927_n803), .Y(_abc_3927_n804_1) );
	NOR2X1 NOR2X1_80 ( .A(_abc_3927_n804_1), .B(_abc_3927_n802), .Y(_abc_3927_n805) );
	AND2X2 AND2X2_53 ( .A(_abc_3927_n799), .B(_abc_3927_n805), .Y(_abc_3927_n806) );
	NAND2X1 NAND2X1_173 ( .A(_abc_3927_n806), .B(_abc_3927_n790_1), .Y(_abc_3927_n807) );
	NAND2X1 NAND2X1_174 ( .A(reg_vv_value_0_), .B(_abc_3927_n480_1), .Y(_abc_3927_n808) );
	NAND2X1 NAND2X1_175 ( .A(_abc_3927_n808), .B(_abc_3927_n766), .Y(_abc_3927_n809_1) );
	NOR2X1 NOR2X1_81 ( .A(_abc_3927_n772), .B(_abc_3927_n809_1), .Y(_abc_3927_n810_1) );
	AND2X2 AND2X2_54 ( .A(_abc_3927_n810_1), .B(_abc_3927_n761), .Y(_abc_3927_n811_1) );
	NAND2X1 NAND2X1_176 ( .A(_abc_3927_n751), .B(_abc_3927_n811_1), .Y(_abc_3927_n812_1) );
	NAND2X1 NAND2X1_177 ( .A(_abc_3927_n812_1), .B(_abc_3927_n807), .Y(_abc_3927_n813_1) );
	NAND2X1 NAND2X1_178 ( .A(_abc_3927_n813_1), .B(_abc_3927_n721), .Y(_abc_3927_n814_1) );
	OR2X2 OR2X2_46 ( .A(_abc_3927_n814_1), .B(_abc_3927_n631), .Y(_abc_3927_n815_1) );
	INVX1 INVX1_33 ( .A(currentaddr_22_), .Y(_abc_3927_n816_1) );
	INVX1 INVX1_34 ( .A(currentaddr_21_), .Y(_abc_3927_n817_1) );
	INVX1 INVX1_35 ( .A(currentaddr_20_), .Y(_abc_3927_n818_1) );
	NOR2X1 NOR2X1_82 ( .A(_abc_3927_n817_1), .B(_abc_3927_n818_1), .Y(_abc_3927_n819_1) );
	INVX1 INVX1_36 ( .A(_abc_3927_n819_1), .Y(_abc_3927_n820_1) );
	NOR2X1 NOR2X1_83 ( .A(_abc_3927_n816_1), .B(_abc_3927_n820_1), .Y(_abc_3927_n821) );
	NAND2X1 NAND2X1_179 ( .A(currentaddr_23_), .B(_abc_3927_n821), .Y(_abc_3927_n822) );
	INVX1 INVX1_37 ( .A(_abc_3927_n822), .Y(_abc_3927_n823) );
	INVX1 INVX1_38 ( .A(currentaddr_19_), .Y(_abc_3927_n824) );
	AND2X2 AND2X2_55 ( .A(currentaddr_17_), .B(currentaddr_16_), .Y(_abc_3927_n825) );
	NAND2X1 NAND2X1_180 ( .A(currentaddr_18_), .B(_abc_3927_n825), .Y(_abc_3927_n826) );
	NOR2X1 NOR2X1_84 ( .A(_abc_3927_n824), .B(_abc_3927_n826), .Y(_abc_3927_n827) );
	INVX1 INVX1_39 ( .A(_abc_3927_n827), .Y(_abc_3927_n828) );
	INVX1 INVX1_40 ( .A(currentaddr_15_), .Y(_abc_3927_n829) );
	INVX1 INVX1_41 ( .A(currentaddr_14_), .Y(_abc_3927_n830) );
	NOR2X1 NOR2X1_85 ( .A(_abc_3927_n829), .B(_abc_3927_n830), .Y(_abc_3927_n831) );
	INVX1 INVX1_42 ( .A(currentaddr_13_), .Y(_abc_3927_n832) );
	INVX2 INVX2_28 ( .A(currentaddr_12_), .Y(_abc_3927_n833) );
	NOR2X1 NOR2X1_86 ( .A(_abc_3927_n832), .B(_abc_3927_n833), .Y(_abc_3927_n834) );
	INVX1 INVX1_43 ( .A(_abc_3927_n834), .Y(_abc_3927_n835) );
	INVX1 INVX1_44 ( .A(currentaddr_11_), .Y(_abc_3927_n836) );
	INVX1 INVX1_45 ( .A(currentaddr_10_), .Y(_abc_3927_n837) );
	NOR2X1 NOR2X1_87 ( .A(_abc_3927_n836), .B(_abc_3927_n837), .Y(_abc_3927_n838) );
	INVX1 INVX1_46 ( .A(currentaddr_6_), .Y(_abc_3927_n839) );
	INVX1 INVX1_47 ( .A(currentaddr_2_), .Y(_abc_3927_n840) );
	NAND2X1 NAND2X1_181 ( .A(currentaddr_1_), .B(currentaddr_0_), .Y(_abc_3927_n841) );
	NOR2X1 NOR2X1_88 ( .A(_abc_3927_n840), .B(_abc_3927_n841), .Y(_abc_3927_n842) );
	AND2X2 AND2X2_56 ( .A(_abc_3927_n842), .B(currentaddr_3_), .Y(_abc_3927_n843) );
	AND2X2 AND2X2_57 ( .A(_abc_3927_n843), .B(currentaddr_4_), .Y(_abc_3927_n844) );
	NAND2X1 NAND2X1_182 ( .A(currentaddr_5_), .B(_abc_3927_n844), .Y(_abc_3927_n845) );
	NOR2X1 NOR2X1_89 ( .A(_abc_3927_n839), .B(_abc_3927_n845), .Y(_abc_3927_n846) );
	NAND2X1 NAND2X1_183 ( .A(currentaddr_7_), .B(_abc_3927_n846), .Y(_abc_3927_n847) );
	INVX1 INVX1_48 ( .A(currentaddr_9_), .Y(_abc_3927_n848) );
	INVX1 INVX1_49 ( .A(currentaddr_8_), .Y(_abc_3927_n849) );
	NOR2X1 NOR2X1_90 ( .A(_abc_3927_n848), .B(_abc_3927_n849), .Y(_abc_3927_n850) );
	INVX1 INVX1_50 ( .A(_abc_3927_n850), .Y(_abc_3927_n851) );
	NOR2X1 NOR2X1_91 ( .A(_abc_3927_n851), .B(_abc_3927_n847), .Y(_abc_3927_n852) );
	NAND2X1 NAND2X1_184 ( .A(_abc_3927_n838), .B(_abc_3927_n852), .Y(_abc_3927_n853) );
	NOR2X1 NOR2X1_92 ( .A(_abc_3927_n835), .B(_abc_3927_n853), .Y(_abc_3927_n854) );
	NAND2X1 NAND2X1_185 ( .A(_abc_3927_n831), .B(_abc_3927_n854), .Y(_abc_3927_n855) );
	NOR2X1 NOR2X1_93 ( .A(_abc_3927_n828), .B(_abc_3927_n855), .Y(_abc_3927_n856) );
	NAND2X1 NAND2X1_186 ( .A(_abc_3927_n823), .B(_abc_3927_n856), .Y(_abc_3927_n857) );
	NOR2X1 NOR2X1_94 ( .A(_abc_3927_n857), .B(_abc_3927_n815_1), .Y(_abc_3927_n858) );
	NAND2X1 NAND2X1_187 ( .A(_abc_3927_n418), .B(_abc_3927_n858), .Y(_abc_3927_n859) );
	XNOR2X1 XNOR2X1_16 ( .A(_abc_3927_n859), .B(_abc_3927_n406), .Y(_abc_3927_n860) );
	NAND2X1 NAND2X1_188 ( .A(_abc_3927_n405), .B(_abc_3927_n860), .Y(_abc_3927_n861) );
	XNOR2X1 XNOR2X1_17 ( .A(currentcol_11_), .B(reg_he_value_11_), .Y(_abc_3927_n862) );
	XNOR2X1 XNOR2X1_18 ( .A(currentcol_10_), .B(reg_he_value_10_), .Y(_abc_3927_n863) );
	NAND2X1 NAND2X1_189 ( .A(_abc_3927_n862), .B(_abc_3927_n863), .Y(_abc_3927_n864) );
	XNOR2X1 XNOR2X1_19 ( .A(currentcol_14_), .B(reg_he_value_14_), .Y(_abc_3927_n865) );
	XNOR2X1 XNOR2X1_20 ( .A(currentcol_15_), .B(reg_he_value_15_), .Y(_abc_3927_n866) );
	NAND2X1 NAND2X1_190 ( .A(_abc_3927_n865), .B(_abc_3927_n866), .Y(_abc_3927_n867) );
	NOR2X1 NOR2X1_95 ( .A(_abc_3927_n864), .B(_abc_3927_n867), .Y(_abc_3927_n868) );
	XNOR2X1 XNOR2X1_21 ( .A(currentcol_0_), .B(reg_he_value_0_), .Y(_abc_3927_n869) );
	XNOR2X1 XNOR2X1_22 ( .A(currentcol_1_), .B(reg_he_value_1_), .Y(_abc_3927_n870) );
	NAND2X1 NAND2X1_191 ( .A(_abc_3927_n869), .B(_abc_3927_n870), .Y(_abc_3927_n871) );
	XNOR2X1 XNOR2X1_23 ( .A(currentcol_4_), .B(reg_he_value_4_), .Y(_abc_3927_n872) );
	XNOR2X1 XNOR2X1_24 ( .A(currentcol_5_), .B(reg_he_value_5_), .Y(_abc_3927_n873) );
	NAND2X1 NAND2X1_192 ( .A(_abc_3927_n872), .B(_abc_3927_n873), .Y(_abc_3927_n874) );
	NOR2X1 NOR2X1_96 ( .A(_abc_3927_n871), .B(_abc_3927_n874), .Y(_abc_3927_n875) );
	NAND2X1 NAND2X1_193 ( .A(_abc_3927_n868), .B(_abc_3927_n875), .Y(_abc_3927_n876) );
	XNOR2X1 XNOR2X1_25 ( .A(currentcol_12_), .B(reg_he_value_12_), .Y(_abc_3927_n877) );
	XNOR2X1 XNOR2X1_26 ( .A(currentcol_13_), .B(reg_he_value_13_), .Y(_abc_3927_n878) );
	NAND2X1 NAND2X1_194 ( .A(_abc_3927_n877), .B(_abc_3927_n878), .Y(_abc_3927_n879) );
	XNOR2X1 XNOR2X1_27 ( .A(currentcol_8_), .B(reg_he_value_8_), .Y(_abc_3927_n880) );
	XNOR2X1 XNOR2X1_28 ( .A(currentcol_9_), .B(reg_he_value_9_), .Y(_abc_3927_n881) );
	NAND2X1 NAND2X1_195 ( .A(_abc_3927_n880), .B(_abc_3927_n881), .Y(_abc_3927_n882) );
	NOR2X1 NOR2X1_97 ( .A(_abc_3927_n879), .B(_abc_3927_n882), .Y(_abc_3927_n883) );
	XNOR2X1 XNOR2X1_29 ( .A(currentcol_3_), .B(reg_he_value_3_), .Y(_abc_3927_n884) );
	XNOR2X1 XNOR2X1_30 ( .A(currentcol_2_), .B(reg_he_value_2_), .Y(_abc_3927_n885) );
	NAND2X1 NAND2X1_196 ( .A(_abc_3927_n884), .B(_abc_3927_n885), .Y(_abc_3927_n886) );
	XNOR2X1 XNOR2X1_31 ( .A(currentcol_7_), .B(reg_he_value_7_), .Y(_abc_3927_n887) );
	XNOR2X1 XNOR2X1_32 ( .A(currentcol_6_), .B(reg_he_value_6_), .Y(_abc_3927_n888) );
	NAND2X1 NAND2X1_197 ( .A(_abc_3927_n887), .B(_abc_3927_n888), .Y(_abc_3927_n889) );
	NOR2X1 NOR2X1_98 ( .A(_abc_3927_n886), .B(_abc_3927_n889), .Y(_abc_3927_n890) );
	NAND2X1 NAND2X1_198 ( .A(_abc_3927_n890), .B(_abc_3927_n883), .Y(_abc_3927_n891) );
	NOR2X1 NOR2X1_99 ( .A(_abc_3927_n876), .B(_abc_3927_n891), .Y(_abc_3927_n892) );
	NOR2X1 NOR2X1_100 ( .A(reg_fh_value_14_), .B(_abc_3927_n405), .Y(_abc_3927_n893) );
	NOR2X1 NOR2X1_101 ( .A(_abc_3927_n892), .B(_abc_3927_n893), .Y(_abc_3927_n894) );
	NAND2X1 NAND2X1_199 ( .A(_abc_3927_n894), .B(_abc_3927_n861), .Y(_abc_3927_n895) );
	AND2X2 AND2X2_58 ( .A(reg_sl_value_1_), .B(currentaddr_1_), .Y(_abc_3927_n896) );
	INVX1 INVX1_51 ( .A(_abc_3927_n896), .Y(_abc_3927_n897) );
	AND2X2 AND2X2_59 ( .A(currentaddr_0_), .B(reg_sl_value_0_), .Y(_abc_3927_n898) );
	NOR2X1 NOR2X1_102 ( .A(reg_sl_value_1_), .B(currentaddr_1_), .Y(_abc_3927_n899) );
	NOR2X1 NOR2X1_103 ( .A(_abc_3927_n899), .B(_abc_3927_n896), .Y(_abc_3927_n900) );
	NAND2X1 NAND2X1_200 ( .A(_abc_3927_n898), .B(_abc_3927_n900), .Y(_abc_3927_n901) );
	NAND2X1 NAND2X1_201 ( .A(_abc_3927_n897), .B(_abc_3927_n901), .Y(_abc_3927_n902) );
	XNOR2X1 XNOR2X1_33 ( .A(currentaddr_3_), .B(reg_sl_value_3_), .Y(_abc_3927_n903) );
	NAND2X1 NAND2X1_202 ( .A(currentaddr_2_), .B(reg_sl_value_2_), .Y(_abc_3927_n904) );
	OR2X2 OR2X2_47 ( .A(currentaddr_2_), .B(reg_sl_value_2_), .Y(_abc_3927_n905) );
	NAND2X1 NAND2X1_203 ( .A(_abc_3927_n904), .B(_abc_3927_n905), .Y(_abc_3927_n906) );
	NOR2X1 NOR2X1_104 ( .A(_abc_3927_n906), .B(_abc_3927_n903), .Y(_abc_3927_n907) );
	NAND2X1 NAND2X1_204 ( .A(_abc_3927_n907), .B(_abc_3927_n902), .Y(_abc_3927_n908) );
	AND2X2 AND2X2_60 ( .A(currentaddr_3_), .B(reg_sl_value_3_), .Y(_abc_3927_n909) );
	NOR2X1 NOR2X1_105 ( .A(_abc_3927_n904), .B(_abc_3927_n903), .Y(_abc_3927_n910) );
	NOR2X1 NOR2X1_106 ( .A(_abc_3927_n909), .B(_abc_3927_n910), .Y(_abc_3927_n911) );
	NAND2X1 NAND2X1_205 ( .A(_abc_3927_n911), .B(_abc_3927_n908), .Y(_abc_3927_n912) );
	NAND2X1 NAND2X1_206 ( .A(reg_sl_value_7_), .B(currentaddr_7_), .Y(_abc_3927_n913) );
	OR2X2 OR2X2_48 ( .A(reg_sl_value_7_), .B(currentaddr_7_), .Y(_abc_3927_n914) );
	AND2X2 AND2X2_61 ( .A(_abc_3927_n914), .B(_abc_3927_n913), .Y(_abc_3927_n915) );
	AND2X2 AND2X2_62 ( .A(currentaddr_6_), .B(reg_sl_value_6_), .Y(_abc_3927_n916) );
	NOR2X1 NOR2X1_107 ( .A(currentaddr_6_), .B(reg_sl_value_6_), .Y(_abc_3927_n917_1) );
	NOR2X1 NOR2X1_108 ( .A(_abc_3927_n917_1), .B(_abc_3927_n916), .Y(_abc_3927_n918) );
	NAND2X1 NAND2X1_207 ( .A(_abc_3927_n918), .B(_abc_3927_n915), .Y(_abc_3927_n919) );
	XOR2X1 XOR2X1_16 ( .A(currentaddr_4_), .B(reg_sl_value_4_), .Y(_abc_3927_n920) );
	NAND2X1 NAND2X1_208 ( .A(currentaddr_5_), .B(reg_sl_value_5_), .Y(_abc_3927_n921) );
	OR2X2 OR2X2_49 ( .A(currentaddr_5_), .B(reg_sl_value_5_), .Y(_abc_3927_n922) );
	AND2X2 AND2X2_63 ( .A(_abc_3927_n922), .B(_abc_3927_n921), .Y(_abc_3927_n923) );
	NAND2X1 NAND2X1_209 ( .A(_abc_3927_n920), .B(_abc_3927_n923), .Y(_abc_3927_n924) );
	NOR2X1 NOR2X1_109 ( .A(_abc_3927_n919), .B(_abc_3927_n924), .Y(_abc_3927_n925) );
	NAND2X1 NAND2X1_210 ( .A(_abc_3927_n925), .B(_abc_3927_n912), .Y(_abc_3927_n926) );
	NAND2X1 NAND2X1_211 ( .A(currentaddr_4_), .B(reg_sl_value_4_), .Y(_abc_3927_n927) );
	NAND2X1 NAND2X1_212 ( .A(_abc_3927_n927), .B(_abc_3927_n921), .Y(_abc_3927_n928) );
	NAND2X1 NAND2X1_213 ( .A(_abc_3927_n922), .B(_abc_3927_n928), .Y(_abc_3927_n929) );
	NOR2X1 NOR2X1_110 ( .A(_abc_3927_n929), .B(_abc_3927_n919), .Y(_abc_3927_n930) );
	NAND2X1 NAND2X1_214 ( .A(_abc_3927_n916), .B(_abc_3927_n914), .Y(_abc_3927_n931) );
	NAND2X1 NAND2X1_215 ( .A(_abc_3927_n913), .B(_abc_3927_n931), .Y(_abc_3927_n932_1) );
	NOR2X1 NOR2X1_111 ( .A(_abc_3927_n932_1), .B(_abc_3927_n930), .Y(_abc_3927_n933_1) );
	NAND2X1 NAND2X1_216 ( .A(_abc_3927_n933_1), .B(_abc_3927_n926), .Y(_abc_3927_n934_1) );
	NAND2X1 NAND2X1_217 ( .A(currentaddr_15_), .B(reg_sl_value_15_), .Y(_abc_3927_n935_1) );
	OR2X2 OR2X2_50 ( .A(currentaddr_15_), .B(reg_sl_value_15_), .Y(_abc_3927_n936_1) );
	AND2X2 AND2X2_64 ( .A(_abc_3927_n936_1), .B(_abc_3927_n935_1), .Y(_abc_3927_n937_1) );
	AND2X2 AND2X2_65 ( .A(currentaddr_14_), .B(reg_sl_value_14_), .Y(_abc_3927_n938_1) );
	NOR2X1 NOR2X1_112 ( .A(currentaddr_14_), .B(reg_sl_value_14_), .Y(_abc_3927_n939_1) );
	NOR2X1 NOR2X1_113 ( .A(_abc_3927_n939_1), .B(_abc_3927_n938_1), .Y(_abc_3927_n940_1) );
	NAND2X1 NAND2X1_218 ( .A(_abc_3927_n940_1), .B(_abc_3927_n937_1), .Y(_abc_3927_n941_1) );
	NAND2X1 NAND2X1_219 ( .A(currentaddr_12_), .B(reg_sl_value_12_), .Y(_abc_3927_n942_1) );
	INVX1 INVX1_52 ( .A(_abc_3927_n942_1), .Y(_abc_3927_n943_1) );
	NOR2X1 NOR2X1_114 ( .A(currentaddr_12_), .B(reg_sl_value_12_), .Y(_abc_3927_n944_1) );
	NOR2X1 NOR2X1_115 ( .A(_abc_3927_n944_1), .B(_abc_3927_n943_1), .Y(_abc_3927_n945_1) );
	INVX1 INVX1_53 ( .A(_abc_3927_n945_1), .Y(_abc_3927_n946_1) );
	NAND2X1 NAND2X1_220 ( .A(currentaddr_13_), .B(reg_sl_value_13_), .Y(_abc_3927_n947) );
	OR2X2 OR2X2_51 ( .A(currentaddr_13_), .B(reg_sl_value_13_), .Y(_abc_3927_n948) );
	NAND2X1 NAND2X1_221 ( .A(_abc_3927_n947), .B(_abc_3927_n948), .Y(_abc_3927_n949) );
	OR2X2 OR2X2_52 ( .A(_abc_3927_n946_1), .B(_abc_3927_n949), .Y(_abc_3927_n950) );
	OR2X2 OR2X2_53 ( .A(_abc_3927_n950), .B(_abc_3927_n941_1), .Y(_abc_3927_n951) );
	AND2X2 AND2X2_66 ( .A(reg_sl_value_11_), .B(currentaddr_11_), .Y(_abc_3927_n952) );
	NOR2X1 NOR2X1_116 ( .A(reg_sl_value_11_), .B(currentaddr_11_), .Y(_abc_3927_n953) );
	NOR2X1 NOR2X1_117 ( .A(_abc_3927_n953), .B(_abc_3927_n952), .Y(_abc_3927_n954) );
	XOR2X1 XOR2X1_17 ( .A(currentaddr_10_), .B(reg_sl_value_10_), .Y(_abc_3927_n955) );
	NAND2X1 NAND2X1_222 ( .A(_abc_3927_n954), .B(_abc_3927_n955), .Y(_abc_3927_n956) );
	NAND2X1 NAND2X1_223 ( .A(currentaddr_9_), .B(reg_sl_value_9_), .Y(_abc_3927_n957) );
	OR2X2 OR2X2_54 ( .A(currentaddr_9_), .B(reg_sl_value_9_), .Y(_abc_3927_n958) );
	NAND2X1 NAND2X1_224 ( .A(_abc_3927_n957), .B(_abc_3927_n958), .Y(_abc_3927_n959) );
	NAND2X1 NAND2X1_225 ( .A(currentaddr_8_), .B(reg_sl_value_8_), .Y(_abc_3927_n960) );
	OR2X2 OR2X2_55 ( .A(currentaddr_8_), .B(reg_sl_value_8_), .Y(_abc_3927_n961) );
	NAND2X1 NAND2X1_226 ( .A(_abc_3927_n960), .B(_abc_3927_n961), .Y(_abc_3927_n962) );
	NOR2X1 NOR2X1_118 ( .A(_abc_3927_n959), .B(_abc_3927_n962), .Y(_abc_3927_n963) );
	INVX1 INVX1_54 ( .A(_abc_3927_n963), .Y(_abc_3927_n964) );
	OR2X2 OR2X2_56 ( .A(_abc_3927_n964), .B(_abc_3927_n956), .Y(_abc_3927_n965) );
	NOR2X1 NOR2X1_119 ( .A(_abc_3927_n965), .B(_abc_3927_n951), .Y(_abc_3927_n966) );
	NAND2X1 NAND2X1_227 ( .A(_abc_3927_n966), .B(_abc_3927_n934_1), .Y(_abc_3927_n967) );
	NOR2X1 NOR2X1_120 ( .A(_abc_3927_n941_1), .B(_abc_3927_n950), .Y(_abc_3927_n968) );
	NAND2X1 NAND2X1_228 ( .A(_abc_3927_n957), .B(_abc_3927_n960), .Y(_abc_3927_n969) );
	NAND2X1 NAND2X1_229 ( .A(_abc_3927_n958), .B(_abc_3927_n969), .Y(_abc_3927_n970) );
	OR2X2 OR2X2_57 ( .A(_abc_3927_n956), .B(_abc_3927_n970), .Y(_abc_3927_n971) );
	NAND2X1 NAND2X1_230 ( .A(currentaddr_10_), .B(reg_sl_value_10_), .Y(_abc_3927_n972_1) );
	NOR2X1 NOR2X1_121 ( .A(_abc_3927_n972_1), .B(_abc_3927_n953), .Y(_abc_3927_n973) );
	NOR2X1 NOR2X1_122 ( .A(_abc_3927_n952), .B(_abc_3927_n973), .Y(_abc_3927_n974) );
	NAND2X1 NAND2X1_231 ( .A(_abc_3927_n974), .B(_abc_3927_n971), .Y(_abc_3927_n975_1) );
	NAND2X1 NAND2X1_232 ( .A(_abc_3927_n975_1), .B(_abc_3927_n968), .Y(_abc_3927_n976) );
	NAND2X1 NAND2X1_233 ( .A(_abc_3927_n942_1), .B(_abc_3927_n947), .Y(_abc_3927_n977) );
	NAND2X1 NAND2X1_234 ( .A(_abc_3927_n948), .B(_abc_3927_n977), .Y(_abc_3927_n978) );
	NOR2X1 NOR2X1_123 ( .A(_abc_3927_n978), .B(_abc_3927_n941_1), .Y(_abc_3927_n979) );
	NAND2X1 NAND2X1_235 ( .A(_abc_3927_n938_1), .B(_abc_3927_n936_1), .Y(_abc_3927_n980) );
	NAND2X1 NAND2X1_236 ( .A(_abc_3927_n935_1), .B(_abc_3927_n980), .Y(_abc_3927_n981_1) );
	NOR2X1 NOR2X1_124 ( .A(_abc_3927_n981_1), .B(_abc_3927_n979), .Y(_abc_3927_n982) );
	AND2X2 AND2X2_67 ( .A(_abc_3927_n976), .B(_abc_3927_n982), .Y(_abc_3927_n983) );
	NAND2X1 NAND2X1_237 ( .A(_abc_3927_n983), .B(_abc_3927_n967), .Y(_abc_3927_n984) );
	AND2X2 AND2X2_68 ( .A(currentaddr_23_), .B(reg_sh_value_7_), .Y(_abc_3927_n985) );
	NOR2X1 NOR2X1_125 ( .A(currentaddr_23_), .B(reg_sh_value_7_), .Y(_abc_3927_n986_1) );
	NOR2X1 NOR2X1_126 ( .A(_abc_3927_n986_1), .B(_abc_3927_n985), .Y(_abc_3927_n987) );
	INVX1 INVX1_55 ( .A(reg_sh_value_6_), .Y(_abc_3927_n988_1) );
	NOR2X1 NOR2X1_127 ( .A(_abc_3927_n816_1), .B(_abc_3927_n988_1), .Y(_abc_3927_n989) );
	NOR2X1 NOR2X1_128 ( .A(currentaddr_22_), .B(reg_sh_value_6_), .Y(_abc_3927_n990) );
	NOR2X1 NOR2X1_129 ( .A(_abc_3927_n990), .B(_abc_3927_n989), .Y(_abc_3927_n991) );
	NAND2X1 NAND2X1_238 ( .A(_abc_3927_n987), .B(_abc_3927_n991), .Y(_abc_3927_n992) );
	NAND2X1 NAND2X1_239 ( .A(reg_sh_value_5_), .B(currentaddr_21_), .Y(_abc_3927_n993_1) );
	NOR2X1 NOR2X1_130 ( .A(reg_sh_value_5_), .B(currentaddr_21_), .Y(_abc_3927_n994) );
	INVX1 INVX1_56 ( .A(_abc_3927_n994), .Y(_abc_3927_n995_1) );
	NAND2X1 NAND2X1_240 ( .A(_abc_3927_n993_1), .B(_abc_3927_n995_1), .Y(_abc_3927_n996) );
	NAND2X1 NAND2X1_241 ( .A(currentaddr_20_), .B(reg_sh_value_4_), .Y(_abc_3927_n997) );
	INVX1 INVX1_57 ( .A(_abc_3927_n997), .Y(_abc_3927_n998) );
	NOR2X1 NOR2X1_131 ( .A(currentaddr_20_), .B(reg_sh_value_4_), .Y(_abc_3927_n999) );
	NOR2X1 NOR2X1_132 ( .A(_abc_3927_n999), .B(_abc_3927_n998), .Y(_abc_3927_n1000_1) );
	INVX1 INVX1_58 ( .A(_abc_3927_n1000_1), .Y(_abc_3927_n1001) );
	NOR2X1 NOR2X1_133 ( .A(_abc_3927_n996), .B(_abc_3927_n1001), .Y(_abc_3927_n1002_1) );
	INVX1 INVX1_59 ( .A(_abc_3927_n1002_1), .Y(_abc_3927_n1003) );
	NOR2X1 NOR2X1_134 ( .A(_abc_3927_n992), .B(_abc_3927_n1003), .Y(_abc_3927_n1004) );
	AND2X2 AND2X2_69 ( .A(currentaddr_19_), .B(reg_sh_value_3_), .Y(_abc_3927_n1005) );
	NOR2X1 NOR2X1_135 ( .A(currentaddr_19_), .B(reg_sh_value_3_), .Y(_abc_3927_n1006) );
	NOR2X1 NOR2X1_136 ( .A(_abc_3927_n1006), .B(_abc_3927_n1005), .Y(_abc_3927_n1007) );
	INVX1 INVX1_60 ( .A(currentaddr_18_), .Y(_abc_3927_n1008) );
	INVX1 INVX1_61 ( .A(reg_sh_value_2_), .Y(_abc_3927_n1009) );
	NOR2X1 NOR2X1_137 ( .A(_abc_3927_n1008), .B(_abc_3927_n1009), .Y(_abc_3927_n1010_1) );
	NOR2X1 NOR2X1_138 ( .A(currentaddr_18_), .B(reg_sh_value_2_), .Y(_abc_3927_n1011_1) );
	NOR2X1 NOR2X1_139 ( .A(_abc_3927_n1011_1), .B(_abc_3927_n1010_1), .Y(_abc_3927_n1012) );
	NAND2X1 NAND2X1_242 ( .A(_abc_3927_n1007), .B(_abc_3927_n1012), .Y(_abc_3927_n1013) );
	INVX1 INVX1_62 ( .A(_abc_3927_n1013), .Y(_abc_3927_n1014) );
	NAND2X1 NAND2X1_243 ( .A(currentaddr_16_), .B(reg_sh_value_0_), .Y(_abc_3927_n1015) );
	INVX1 INVX1_63 ( .A(_abc_3927_n1015), .Y(_abc_3927_n1016) );
	NOR2X1 NOR2X1_140 ( .A(currentaddr_16_), .B(reg_sh_value_0_), .Y(_abc_3927_n1017) );
	NOR2X1 NOR2X1_141 ( .A(_abc_3927_n1017), .B(_abc_3927_n1016), .Y(_abc_3927_n1018) );
	INVX1 INVX1_64 ( .A(_abc_3927_n1018), .Y(_abc_3927_n1019) );
	NAND2X1 NAND2X1_244 ( .A(reg_sh_value_1_), .B(currentaddr_17_), .Y(_abc_3927_n1020) );
	NOR2X1 NOR2X1_142 ( .A(reg_sh_value_1_), .B(currentaddr_17_), .Y(_abc_3927_n1021) );
	INVX1 INVX1_65 ( .A(_abc_3927_n1021), .Y(_abc_3927_n1022) );
	NAND2X1 NAND2X1_245 ( .A(_abc_3927_n1020), .B(_abc_3927_n1022), .Y(_abc_3927_n1023) );
	NOR2X1 NOR2X1_143 ( .A(_abc_3927_n1023), .B(_abc_3927_n1019), .Y(_abc_3927_n1024_1) );
	NAND2X1 NAND2X1_246 ( .A(_abc_3927_n1024_1), .B(_abc_3927_n1014), .Y(_abc_3927_n1025) );
	INVX1 INVX1_66 ( .A(_abc_3927_n1025), .Y(_abc_3927_n1026) );
	AND2X2 AND2X2_70 ( .A(_abc_3927_n1004), .B(_abc_3927_n1026), .Y(_abc_3927_n1027) );
	NAND2X1 NAND2X1_247 ( .A(_abc_3927_n1027), .B(_abc_3927_n984), .Y(_abc_3927_n1028_1) );
	NAND2X1 NAND2X1_248 ( .A(_abc_3927_n993_1), .B(_abc_3927_n997), .Y(_abc_3927_n1029) );
	NAND2X1 NAND2X1_249 ( .A(_abc_3927_n1029), .B(_abc_3927_n995_1), .Y(_abc_3927_n1030) );
	NOR2X1 NOR2X1_144 ( .A(_abc_3927_n1030), .B(_abc_3927_n992), .Y(_abc_3927_n1031) );
	NAND2X1 NAND2X1_250 ( .A(_abc_3927_n1015), .B(_abc_3927_n1020), .Y(_abc_3927_n1032) );
	NAND2X1 NAND2X1_251 ( .A(_abc_3927_n1032), .B(_abc_3927_n1022), .Y(_abc_3927_n1033) );
	OR2X2 OR2X2_58 ( .A(_abc_3927_n1013), .B(_abc_3927_n1033), .Y(_abc_3927_n1034) );
	INVX1 INVX1_67 ( .A(_abc_3927_n1010_1), .Y(_abc_3927_n1035) );
	NOR2X1 NOR2X1_145 ( .A(_abc_3927_n1006), .B(_abc_3927_n1035), .Y(_abc_3927_n1036_1) );
	NOR2X1 NOR2X1_146 ( .A(_abc_3927_n1005), .B(_abc_3927_n1036_1), .Y(_abc_3927_n1037_1) );
	NAND2X1 NAND2X1_252 ( .A(_abc_3927_n1037_1), .B(_abc_3927_n1034), .Y(_abc_3927_n1038) );
	NAND2X1 NAND2X1_253 ( .A(_abc_3927_n1038), .B(_abc_3927_n1004), .Y(_abc_3927_n1039) );
	INVX1 INVX1_68 ( .A(_abc_3927_n989), .Y(_abc_3927_n1040) );
	NOR2X1 NOR2X1_147 ( .A(_abc_3927_n986_1), .B(_abc_3927_n1040), .Y(_abc_3927_n1041) );
	NOR2X1 NOR2X1_148 ( .A(_abc_3927_n985), .B(_abc_3927_n1041), .Y(_abc_3927_n1042) );
	NAND2X1 NAND2X1_254 ( .A(_abc_3927_n1042), .B(_abc_3927_n1039), .Y(_abc_3927_n1043) );
	NOR2X1 NOR2X1_149 ( .A(_abc_3927_n1031), .B(_abc_3927_n1043), .Y(_abc_3927_n1044) );
	NAND2X1 NAND2X1_255 ( .A(_abc_3927_n1044), .B(_abc_3927_n1028_1), .Y(_abc_3927_n1045) );
	AND2X2 AND2X2_71 ( .A(currentaddr_27_), .B(reg_sh_value_11_), .Y(_abc_3927_n1046) );
	NOR2X1 NOR2X1_150 ( .A(currentaddr_27_), .B(reg_sh_value_11_), .Y(_abc_3927_n1047_1) );
	NOR2X1 NOR2X1_151 ( .A(_abc_3927_n1047_1), .B(_abc_3927_n1046), .Y(_abc_3927_n1048) );
	INVX1 INVX1_69 ( .A(reg_sh_value_10_), .Y(_abc_3927_n1049) );
	NOR2X1 NOR2X1_152 ( .A(_abc_3927_n414), .B(_abc_3927_n1049), .Y(_abc_3927_n1050) );
	NOR2X1 NOR2X1_153 ( .A(currentaddr_26_), .B(reg_sh_value_10_), .Y(_abc_3927_n1051) );
	NOR2X1 NOR2X1_154 ( .A(_abc_3927_n1051), .B(_abc_3927_n1050), .Y(_abc_3927_n1052) );
	NAND2X1 NAND2X1_256 ( .A(_abc_3927_n1048), .B(_abc_3927_n1052), .Y(_abc_3927_n1053) );
	AND2X2 AND2X2_72 ( .A(reg_sh_value_9_), .B(currentaddr_25_), .Y(_abc_3927_n1054) );
	NOR2X1 NOR2X1_155 ( .A(reg_sh_value_9_), .B(currentaddr_25_), .Y(_abc_3927_n1055) );
	NOR2X1 NOR2X1_156 ( .A(_abc_3927_n1055), .B(_abc_3927_n1054), .Y(_abc_3927_n1056) );
	INVX1 INVX1_70 ( .A(reg_sh_value_8_), .Y(_abc_3927_n1057) );
	NOR2X1 NOR2X1_157 ( .A(_abc_3927_n411), .B(_abc_3927_n1057), .Y(_abc_3927_n1058_1) );
	NOR2X1 NOR2X1_158 ( .A(currentaddr_24_), .B(reg_sh_value_8_), .Y(_abc_3927_n1059) );
	NOR2X1 NOR2X1_159 ( .A(_abc_3927_n1059), .B(_abc_3927_n1058_1), .Y(_abc_3927_n1060) );
	NAND2X1 NAND2X1_257 ( .A(_abc_3927_n1056), .B(_abc_3927_n1060), .Y(_abc_3927_n1061) );
	NOR2X1 NOR2X1_160 ( .A(_abc_3927_n1053), .B(_abc_3927_n1061), .Y(_abc_3927_n1062_1) );
	NAND2X1 NAND2X1_258 ( .A(_abc_3927_n1062_1), .B(_abc_3927_n1045), .Y(_abc_3927_n1063) );
	NOR2X1 NOR2X1_161 ( .A(_abc_3927_n1054), .B(_abc_3927_n1058_1), .Y(_abc_3927_n1064) );
	OR2X2 OR2X2_59 ( .A(_abc_3927_n1064), .B(_abc_3927_n1055), .Y(_abc_3927_n1065_1) );
	NOR2X1 NOR2X1_162 ( .A(_abc_3927_n1053), .B(_abc_3927_n1065_1), .Y(_abc_3927_n1066_1) );
	INVX1 INVX1_71 ( .A(_abc_3927_n1050), .Y(_abc_3927_n1067) );
	NOR2X1 NOR2X1_163 ( .A(_abc_3927_n1047_1), .B(_abc_3927_n1067), .Y(_abc_3927_n1068_1) );
	OR2X2 OR2X2_60 ( .A(_abc_3927_n1068_1), .B(_abc_3927_n1046), .Y(_abc_3927_n1069) );
	NOR2X1 NOR2X1_164 ( .A(_abc_3927_n1069), .B(_abc_3927_n1066_1), .Y(_abc_3927_n1070_1) );
	NAND2X1 NAND2X1_259 ( .A(_abc_3927_n1070_1), .B(_abc_3927_n1063), .Y(_abc_3927_n1071) );
	AND2X2 AND2X2_73 ( .A(currentaddr_29_), .B(reg_sh_value_13_), .Y(_abc_3927_n1072_1) );
	NOR2X1 NOR2X1_165 ( .A(currentaddr_29_), .B(reg_sh_value_13_), .Y(_abc_3927_n1073) );
	OR2X2 OR2X2_61 ( .A(_abc_3927_n1072_1), .B(_abc_3927_n1073), .Y(_abc_3927_n1074_1) );
	INVX1 INVX1_72 ( .A(reg_sh_value_12_), .Y(_abc_3927_n1075) );
	NOR2X1 NOR2X1_166 ( .A(_abc_3927_n407), .B(_abc_3927_n1075), .Y(_abc_3927_n1076_1) );
	NOR2X1 NOR2X1_167 ( .A(currentaddr_28_), .B(reg_sh_value_12_), .Y(_abc_3927_n1077) );
	NOR2X1 NOR2X1_168 ( .A(_abc_3927_n1077), .B(_abc_3927_n1076_1), .Y(_abc_3927_n1078_1) );
	INVX1 INVX1_73 ( .A(_abc_3927_n1078_1), .Y(_abc_3927_n1079) );
	NOR2X1 NOR2X1_169 ( .A(_abc_3927_n1074_1), .B(_abc_3927_n1079), .Y(_abc_3927_n1080_1) );
	NAND2X1 NAND2X1_260 ( .A(_abc_3927_n1080_1), .B(_abc_3927_n1071), .Y(_abc_3927_n1081) );
	INVX1 INVX1_74 ( .A(_abc_3927_n1076_1), .Y(_abc_3927_n1082_1) );
	NOR2X1 NOR2X1_170 ( .A(_abc_3927_n1073), .B(_abc_3927_n1082_1), .Y(_abc_3927_n1083) );
	NOR2X1 NOR2X1_171 ( .A(_abc_3927_n1072_1), .B(_abc_3927_n1083), .Y(_abc_3927_n1084_1) );
	NAND2X1 NAND2X1_261 ( .A(_abc_3927_n1084_1), .B(_abc_3927_n1081), .Y(_abc_3927_n1085) );
	XOR2X1 XOR2X1_18 ( .A(currentaddr_30_), .B(reg_sh_value_14_), .Y(_abc_3927_n1086_1) );
	NAND2X1 NAND2X1_262 ( .A(_abc_3927_n1086_1), .B(_abc_3927_n1085), .Y(_abc_3927_n1087) );
	INVX4 INVX4_2 ( .A(_abc_3927_n892), .Y(_abc_3927_n1088_1) );
	NOR2X1 NOR2X1_172 ( .A(_abc_3927_n1086_1), .B(_abc_3927_n1085), .Y(_abc_3927_n1089) );
	NOR2X1 NOR2X1_173 ( .A(_abc_3927_n1088_1), .B(_abc_3927_n1089), .Y(_abc_3927_n1090_1) );
	NAND2X1 NAND2X1_263 ( .A(_abc_3927_n1087), .B(_abc_3927_n1090_1), .Y(_abc_3927_n1091) );
	NAND2X1 NAND2X1_264 ( .A(_abc_3927_n1091), .B(_abc_3927_n895), .Y(_abc_3927_n1092_1) );
	AND2X2 AND2X2_74 ( .A(_abc_3927_n1092_1), .B(_abc_3927_n365), .Y(currentaddr_30__FF_INPUT) );
	NOR2X1 NOR2X1_174 ( .A(_abc_3927_n631), .B(_abc_3927_n814_1), .Y(_abc_3927_n1094_1) );
	NOR2X1 NOR2X1_175 ( .A(_abc_3927_n408), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1095) );
	NOR2X1 NOR2X1_176 ( .A(_abc_3927_n828), .B(_abc_3927_n822), .Y(_abc_3927_n1096_1) );
	INVX1 INVX1_75 ( .A(_abc_3927_n831), .Y(_abc_3927_n1097) );
	NOR2X1 NOR2X1_177 ( .A(_abc_3927_n835), .B(_abc_3927_n1097), .Y(_abc_3927_n1098_1) );
	INVX1 INVX1_76 ( .A(_abc_3927_n838), .Y(_abc_3927_n1099) );
	NOR2X1 NOR2X1_178 ( .A(_abc_3927_n851), .B(_abc_3927_n1099), .Y(_abc_3927_n1100_1) );
	NAND2X1 NAND2X1_265 ( .A(_abc_3927_n1098_1), .B(_abc_3927_n1100_1), .Y(_abc_3927_n1101) );
	NAND2X1 NAND2X1_266 ( .A(currentaddr_5_), .B(currentaddr_4_), .Y(_abc_3927_n1102_1) );
	NAND2X1 NAND2X1_267 ( .A(currentaddr_7_), .B(currentaddr_6_), .Y(_abc_3927_n1103) );
	NOR2X1 NOR2X1_179 ( .A(_abc_3927_n1102_1), .B(_abc_3927_n1103), .Y(_abc_3927_n1104_1) );
	NAND2X1 NAND2X1_268 ( .A(_abc_3927_n1104_1), .B(_abc_3927_n843), .Y(_abc_3927_n1105) );
	NOR2X1 NOR2X1_180 ( .A(_abc_3927_n1105), .B(_abc_3927_n1101), .Y(_abc_3927_n1106_1) );
	NAND2X1 NAND2X1_269 ( .A(_abc_3927_n1096_1), .B(_abc_3927_n1106_1), .Y(_abc_3927_n1107) );
	NOR2X1 NOR2X1_181 ( .A(_abc_3927_n416), .B(_abc_3927_n1107), .Y(_abc_3927_n1108_1) );
	NAND2X1 NAND2X1_270 ( .A(currentaddr_28_), .B(_abc_3927_n1108_1), .Y(_abc_3927_n1109) );
	XNOR2X1 XNOR2X1_34 ( .A(_abc_3927_n1109), .B(currentaddr_29_), .Y(_abc_3927_n1110_1) );
	AND2X2 AND2X2_75 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1110_1), .Y(_abc_3927_n1111) );
	NOR2X1 NOR2X1_182 ( .A(_abc_3927_n1095), .B(_abc_3927_n1111), .Y(_abc_3927_n1112_1) );
	NAND2X1 NAND2X1_271 ( .A(_abc_3927_n405), .B(_abc_3927_n1112_1), .Y(_abc_3927_n1113) );
	NOR2X1 NOR2X1_183 ( .A(reg_fh_value_13_), .B(_abc_3927_n405), .Y(_abc_3927_n1114_1) );
	NOR2X1 NOR2X1_184 ( .A(_abc_3927_n892), .B(_abc_3927_n1114_1), .Y(_abc_3927_n1115) );
	NAND2X1 NAND2X1_272 ( .A(_abc_3927_n1115), .B(_abc_3927_n1113), .Y(_abc_3927_n1116_1) );
	NAND2X1 NAND2X1_273 ( .A(_abc_3927_n1078_1), .B(_abc_3927_n1071), .Y(_abc_3927_n1117) );
	NAND2X1 NAND2X1_274 ( .A(_abc_3927_n1082_1), .B(_abc_3927_n1117), .Y(_abc_3927_n1118_1) );
	XNOR2X1 XNOR2X1_35 ( .A(_abc_3927_n1118_1), .B(_abc_3927_n1074_1), .Y(_abc_3927_n1119) );
	NAND2X1 NAND2X1_275 ( .A(_abc_3927_n892), .B(_abc_3927_n1119), .Y(_abc_3927_n1120_1) );
	NAND2X1 NAND2X1_276 ( .A(_abc_3927_n1116_1), .B(_abc_3927_n1120_1), .Y(_abc_3927_n1121) );
	AND2X2 AND2X2_76 ( .A(_abc_3927_n1121), .B(_abc_3927_n365), .Y(currentaddr_29__FF_INPUT) );
	NAND2X1 NAND2X1_277 ( .A(_abc_3927_n417), .B(_abc_3927_n858), .Y(_abc_3927_n1123) );
	XNOR2X1 XNOR2X1_36 ( .A(_abc_3927_n1123), .B(_abc_3927_n407), .Y(_abc_3927_n1124_1) );
	NAND2X1 NAND2X1_278 ( .A(_abc_3927_n405), .B(_abc_3927_n1124_1), .Y(_abc_3927_n1125) );
	NOR2X1 NOR2X1_185 ( .A(reg_fh_value_12_), .B(_abc_3927_n405), .Y(_abc_3927_n1126_1) );
	NOR2X1 NOR2X1_186 ( .A(_abc_3927_n892), .B(_abc_3927_n1126_1), .Y(_abc_3927_n1127) );
	NAND2X1 NAND2X1_279 ( .A(_abc_3927_n1127), .B(_abc_3927_n1125), .Y(_abc_3927_n1128_1) );
	XNOR2X1 XNOR2X1_37 ( .A(_abc_3927_n1071), .B(_abc_3927_n1079), .Y(_abc_3927_n1129) );
	NAND2X1 NAND2X1_280 ( .A(_abc_3927_n892), .B(_abc_3927_n1129), .Y(_abc_3927_n1130_1) );
	NAND2X1 NAND2X1_281 ( .A(_abc_3927_n1130_1), .B(_abc_3927_n1128_1), .Y(_abc_3927_n1131) );
	AND2X2 AND2X2_77 ( .A(_abc_3927_n1131), .B(_abc_3927_n365), .Y(currentaddr_28__FF_INPUT) );
	NOR2X1 NOR2X1_187 ( .A(_abc_3927_n413), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1133) );
	INVX1 INVX1_77 ( .A(_abc_3927_n412), .Y(_abc_3927_n1134_1) );
	NOR2X1 NOR2X1_188 ( .A(_abc_3927_n1134_1), .B(_abc_3927_n1107), .Y(_abc_3927_n1135) );
	NAND2X1 NAND2X1_282 ( .A(currentaddr_26_), .B(_abc_3927_n1135), .Y(_abc_3927_n1136_1) );
	XNOR2X1 XNOR2X1_38 ( .A(_abc_3927_n1136_1), .B(currentaddr_27_), .Y(_abc_3927_n1137) );
	AND2X2 AND2X2_78 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1137), .Y(_abc_3927_n1138_1) );
	NOR2X1 NOR2X1_189 ( .A(_abc_3927_n1133), .B(_abc_3927_n1138_1), .Y(_abc_3927_n1139) );
	NAND2X1 NAND2X1_283 ( .A(_abc_3927_n405), .B(_abc_3927_n1139), .Y(_abc_3927_n1140_1) );
	NOR2X1 NOR2X1_190 ( .A(reg_fh_value_11_), .B(_abc_3927_n405), .Y(_abc_3927_n1141) );
	NOR2X1 NOR2X1_191 ( .A(_abc_3927_n892), .B(_abc_3927_n1141), .Y(_abc_3927_n1142_1) );
	NAND2X1 NAND2X1_284 ( .A(_abc_3927_n1142_1), .B(_abc_3927_n1140_1), .Y(_abc_3927_n1143) );
	NAND2X1 NAND2X1_285 ( .A(_abc_3927_n1060), .B(_abc_3927_n1045), .Y(_abc_3927_n1144_1) );
	AND2X2 AND2X2_79 ( .A(_abc_3927_n1144_1), .B(_abc_3927_n1064), .Y(_abc_3927_n1145) );
	NOR2X1 NOR2X1_192 ( .A(_abc_3927_n1055), .B(_abc_3927_n1145), .Y(_abc_3927_n1146_1) );
	NAND2X1 NAND2X1_286 ( .A(_abc_3927_n1052), .B(_abc_3927_n1146_1), .Y(_abc_3927_n1147) );
	NAND2X1 NAND2X1_287 ( .A(_abc_3927_n1067), .B(_abc_3927_n1147), .Y(_abc_3927_n1148_1) );
	XOR2X1 XOR2X1_19 ( .A(_abc_3927_n1148_1), .B(_abc_3927_n1048), .Y(_abc_3927_n1149) );
	NAND2X1 NAND2X1_288 ( .A(_abc_3927_n892), .B(_abc_3927_n1149), .Y(_abc_3927_n1150_1) );
	NAND2X1 NAND2X1_289 ( .A(_abc_3927_n1143), .B(_abc_3927_n1150_1), .Y(_abc_3927_n1151) );
	AND2X2 AND2X2_80 ( .A(_abc_3927_n1151), .B(_abc_3927_n365), .Y(currentaddr_27__FF_INPUT) );
	NAND2X1 NAND2X1_290 ( .A(_abc_3927_n412), .B(_abc_3927_n858), .Y(_abc_3927_n1153) );
	XNOR2X1 XNOR2X1_39 ( .A(_abc_3927_n1153), .B(_abc_3927_n414), .Y(_abc_3927_n1154_1) );
	NAND2X1 NAND2X1_291 ( .A(_abc_3927_n405), .B(_abc_3927_n1154_1), .Y(_abc_3927_n1155) );
	NOR2X1 NOR2X1_193 ( .A(reg_fh_value_10_), .B(_abc_3927_n405), .Y(_abc_3927_n1156_1) );
	NOR2X1 NOR2X1_194 ( .A(_abc_3927_n892), .B(_abc_3927_n1156_1), .Y(_abc_3927_n1157) );
	NAND2X1 NAND2X1_292 ( .A(_abc_3927_n1157), .B(_abc_3927_n1155), .Y(_abc_3927_n1158_1) );
	NOR2X1 NOR2X1_195 ( .A(_abc_3927_n1052), .B(_abc_3927_n1146_1), .Y(_abc_3927_n1159) );
	NAND2X1 NAND2X1_293 ( .A(_abc_3927_n892), .B(_abc_3927_n1147), .Y(_abc_3927_n1160_1) );
	OR2X2 OR2X2_62 ( .A(_abc_3927_n1160_1), .B(_abc_3927_n1159), .Y(_abc_3927_n1161) );
	NAND2X1 NAND2X1_294 ( .A(_abc_3927_n1161), .B(_abc_3927_n1158_1), .Y(_abc_3927_n1162_1) );
	AND2X2 AND2X2_81 ( .A(_abc_3927_n1162_1), .B(_abc_3927_n365), .Y(currentaddr_26__FF_INPUT) );
	NAND2X1 NAND2X1_295 ( .A(currentaddr_24_), .B(_abc_3927_n858), .Y(_abc_3927_n1164_1) );
	XNOR2X1 XNOR2X1_40 ( .A(_abc_3927_n1164_1), .B(_abc_3927_n410), .Y(_abc_3927_n1165) );
	NAND2X1 NAND2X1_296 ( .A(_abc_3927_n405), .B(_abc_3927_n1165), .Y(_abc_3927_n1166_1) );
	NOR2X1 NOR2X1_196 ( .A(reg_fh_value_9_), .B(_abc_3927_n405), .Y(_abc_3927_n1167) );
	NOR2X1 NOR2X1_197 ( .A(_abc_3927_n892), .B(_abc_3927_n1167), .Y(_abc_3927_n1168_1) );
	NAND2X1 NAND2X1_297 ( .A(_abc_3927_n1168_1), .B(_abc_3927_n1166_1), .Y(_abc_3927_n1169) );
	INVX1 INVX1_78 ( .A(_abc_3927_n1058_1), .Y(_abc_3927_n1170_1) );
	NAND2X1 NAND2X1_298 ( .A(_abc_3927_n1170_1), .B(_abc_3927_n1144_1), .Y(_abc_3927_n1171) );
	XOR2X1 XOR2X1_20 ( .A(_abc_3927_n1171), .B(_abc_3927_n1056), .Y(_abc_3927_n1172_1) );
	NAND2X1 NAND2X1_299 ( .A(_abc_3927_n892), .B(_abc_3927_n1172_1), .Y(_abc_3927_n1173) );
	NAND2X1 NAND2X1_300 ( .A(_abc_3927_n1173), .B(_abc_3927_n1169), .Y(_abc_3927_n1174_1) );
	AND2X2 AND2X2_82 ( .A(_abc_3927_n1174_1), .B(_abc_3927_n365), .Y(currentaddr_25__FF_INPUT) );
	NOR2X1 NOR2X1_198 ( .A(_abc_3927_n835), .B(_abc_3927_n1099), .Y(_abc_3927_n1176_1) );
	NAND2X1 NAND2X1_301 ( .A(_abc_3927_n850), .B(_abc_3927_n1176_1), .Y(_abc_3927_n1177) );
	NOR2X1 NOR2X1_199 ( .A(_abc_3927_n1177), .B(_abc_3927_n847), .Y(_abc_3927_n1178_1) );
	INVX1 INVX1_79 ( .A(_abc_3927_n1178_1), .Y(_abc_3927_n1179) );
	NOR2X1 NOR2X1_200 ( .A(_abc_3927_n826), .B(_abc_3927_n1097), .Y(_abc_3927_n1180_1) );
	NAND2X1 NAND2X1_302 ( .A(currentaddr_19_), .B(_abc_3927_n1180_1), .Y(_abc_3927_n1181) );
	NOR2X1 NOR2X1_201 ( .A(_abc_3927_n1181), .B(_abc_3927_n1179), .Y(_abc_3927_n1182_1) );
	NAND2X1 NAND2X1_303 ( .A(_abc_3927_n1182_1), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1183) );
	INVX1 INVX1_80 ( .A(_abc_3927_n1183), .Y(_abc_3927_n1184_1) );
	NAND2X1 NAND2X1_304 ( .A(_abc_3927_n823), .B(_abc_3927_n1184_1), .Y(_abc_3927_n1185) );
	NAND2X1 NAND2X1_305 ( .A(_abc_3927_n411), .B(_abc_3927_n1185), .Y(_abc_3927_n1186_1) );
	NAND2X1 NAND2X1_306 ( .A(_abc_3927_n1164_1), .B(_abc_3927_n1186_1), .Y(_abc_3927_n1187) );
	NAND2X1 NAND2X1_307 ( .A(_abc_3927_n405), .B(_abc_3927_n1187), .Y(_abc_3927_n1188) );
	NOR2X1 NOR2X1_202 ( .A(reg_fh_value_8_), .B(_abc_3927_n405), .Y(_abc_3927_n1189) );
	NOR2X1 NOR2X1_203 ( .A(_abc_3927_n892), .B(_abc_3927_n1189), .Y(_abc_3927_n1190) );
	NAND2X1 NAND2X1_308 ( .A(_abc_3927_n1190), .B(_abc_3927_n1188), .Y(_abc_3927_n1191) );
	XOR2X1 XOR2X1_21 ( .A(_abc_3927_n1045), .B(_abc_3927_n1060), .Y(_abc_3927_n1192) );
	NAND2X1 NAND2X1_309 ( .A(_abc_3927_n892), .B(_abc_3927_n1192), .Y(_abc_3927_n1193) );
	NAND2X1 NAND2X1_310 ( .A(_abc_3927_n1193), .B(_abc_3927_n1191), .Y(_abc_3927_n1194) );
	AND2X2 AND2X2_83 ( .A(_abc_3927_n1194), .B(_abc_3927_n365), .Y(currentaddr_24__FF_INPUT) );
	INVX1 INVX1_81 ( .A(currentaddr_23_), .Y(_abc_3927_n1196) );
	NAND2X1 NAND2X1_311 ( .A(_abc_3927_n821), .B(_abc_3927_n1184_1), .Y(_abc_3927_n1197) );
	NAND2X1 NAND2X1_312 ( .A(_abc_3927_n1196), .B(_abc_3927_n1197), .Y(_abc_3927_n1198) );
	NAND2X1 NAND2X1_313 ( .A(_abc_3927_n1185), .B(_abc_3927_n1198), .Y(_abc_3927_n1199) );
	NAND2X1 NAND2X1_314 ( .A(_abc_3927_n405), .B(_abc_3927_n1199), .Y(_abc_3927_n1200) );
	NOR2X1 NOR2X1_204 ( .A(reg_fh_value_7_), .B(_abc_3927_n405), .Y(_abc_3927_n1201) );
	NOR2X1 NOR2X1_205 ( .A(_abc_3927_n892), .B(_abc_3927_n1201), .Y(_abc_3927_n1202) );
	NAND2X1 NAND2X1_315 ( .A(_abc_3927_n1202), .B(_abc_3927_n1200), .Y(_abc_3927_n1203) );
	INVX1 INVX1_82 ( .A(_abc_3927_n1038), .Y(_abc_3927_n1204) );
	NAND2X1 NAND2X1_316 ( .A(_abc_3927_n1026), .B(_abc_3927_n984), .Y(_abc_3927_n1205) );
	NAND2X1 NAND2X1_317 ( .A(_abc_3927_n1204), .B(_abc_3927_n1205), .Y(_abc_3927_n1206) );
	NAND2X1 NAND2X1_318 ( .A(_abc_3927_n1002_1), .B(_abc_3927_n1206), .Y(_abc_3927_n1207) );
	NAND2X1 NAND2X1_319 ( .A(_abc_3927_n1030), .B(_abc_3927_n1207), .Y(_abc_3927_n1208) );
	NAND2X1 NAND2X1_320 ( .A(_abc_3927_n991), .B(_abc_3927_n1208), .Y(_abc_3927_n1209) );
	NAND2X1 NAND2X1_321 ( .A(_abc_3927_n1040), .B(_abc_3927_n1209), .Y(_abc_3927_n1210) );
	XOR2X1 XOR2X1_22 ( .A(_abc_3927_n1210), .B(_abc_3927_n987), .Y(_abc_3927_n1211) );
	NAND2X1 NAND2X1_322 ( .A(_abc_3927_n892), .B(_abc_3927_n1211), .Y(_abc_3927_n1212) );
	NAND2X1 NAND2X1_323 ( .A(_abc_3927_n1212), .B(_abc_3927_n1203), .Y(_abc_3927_n1213) );
	AND2X2 AND2X2_84 ( .A(_abc_3927_n1213), .B(_abc_3927_n365), .Y(currentaddr_23__FF_INPUT) );
	NAND2X1 NAND2X1_324 ( .A(_abc_3927_n819_1), .B(_abc_3927_n1184_1), .Y(_abc_3927_n1215) );
	NAND2X1 NAND2X1_325 ( .A(_abc_3927_n816_1), .B(_abc_3927_n1215), .Y(_abc_3927_n1216) );
	NAND2X1 NAND2X1_326 ( .A(_abc_3927_n1197), .B(_abc_3927_n1216), .Y(_abc_3927_n1217) );
	NAND2X1 NAND2X1_327 ( .A(_abc_3927_n405), .B(_abc_3927_n1217), .Y(_abc_3927_n1218) );
	NOR2X1 NOR2X1_206 ( .A(reg_fh_value_6_), .B(_abc_3927_n405), .Y(_abc_3927_n1219) );
	NOR2X1 NOR2X1_207 ( .A(_abc_3927_n892), .B(_abc_3927_n1219), .Y(_abc_3927_n1220) );
	NAND2X1 NAND2X1_328 ( .A(_abc_3927_n1220), .B(_abc_3927_n1218), .Y(_abc_3927_n1221) );
	NOR2X1 NOR2X1_208 ( .A(_abc_3927_n991), .B(_abc_3927_n1208), .Y(_abc_3927_n1222_1) );
	NAND2X1 NAND2X1_329 ( .A(_abc_3927_n892), .B(_abc_3927_n1209), .Y(_abc_3927_n1223) );
	OR2X2 OR2X2_63 ( .A(_abc_3927_n1223), .B(_abc_3927_n1222_1), .Y(_abc_3927_n1224) );
	NAND2X1 NAND2X1_330 ( .A(_abc_3927_n1224), .B(_abc_3927_n1221), .Y(_abc_3927_n1225_1) );
	AND2X2 AND2X2_85 ( .A(_abc_3927_n1225_1), .B(_abc_3927_n365), .Y(currentaddr_22__FF_INPUT) );
	NAND2X1 NAND2X1_331 ( .A(currentaddr_20_), .B(_abc_3927_n1184_1), .Y(_abc_3927_n1227_1) );
	NAND2X1 NAND2X1_332 ( .A(_abc_3927_n817_1), .B(_abc_3927_n1227_1), .Y(_abc_3927_n1228) );
	NAND2X1 NAND2X1_333 ( .A(_abc_3927_n1215), .B(_abc_3927_n1228), .Y(_abc_3927_n1229_1) );
	NAND2X1 NAND2X1_334 ( .A(_abc_3927_n405), .B(_abc_3927_n1229_1), .Y(_abc_3927_n1230) );
	NOR2X1 NOR2X1_209 ( .A(reg_fh_value_5_), .B(_abc_3927_n405), .Y(_abc_3927_n1231_1) );
	NOR2X1 NOR2X1_210 ( .A(_abc_3927_n892), .B(_abc_3927_n1231_1), .Y(_abc_3927_n1232) );
	NAND2X1 NAND2X1_335 ( .A(_abc_3927_n1232), .B(_abc_3927_n1230), .Y(_abc_3927_n1233_1) );
	NAND2X1 NAND2X1_336 ( .A(_abc_3927_n1000_1), .B(_abc_3927_n1206), .Y(_abc_3927_n1234) );
	NAND2X1 NAND2X1_337 ( .A(_abc_3927_n997), .B(_abc_3927_n1234), .Y(_abc_3927_n1235_1) );
	XNOR2X1 XNOR2X1_41 ( .A(_abc_3927_n1235_1), .B(_abc_3927_n996), .Y(_abc_3927_n1236) );
	NAND2X1 NAND2X1_338 ( .A(_abc_3927_n892), .B(_abc_3927_n1236), .Y(_abc_3927_n1237_1) );
	NAND2X1 NAND2X1_339 ( .A(_abc_3927_n1237_1), .B(_abc_3927_n1233_1), .Y(_abc_3927_n1238) );
	AND2X2 AND2X2_86 ( .A(_abc_3927_n1238), .B(_abc_3927_n365), .Y(currentaddr_21__FF_INPUT) );
	NAND2X1 NAND2X1_340 ( .A(_abc_3927_n818_1), .B(_abc_3927_n1183), .Y(_abc_3927_n1240) );
	NAND2X1 NAND2X1_341 ( .A(_abc_3927_n1240), .B(_abc_3927_n1227_1), .Y(_abc_3927_n1241_1) );
	NAND2X1 NAND2X1_342 ( .A(_abc_3927_n405), .B(_abc_3927_n1241_1), .Y(_abc_3927_n1242) );
	NOR2X1 NOR2X1_211 ( .A(reg_fh_value_4_), .B(_abc_3927_n405), .Y(_abc_3927_n1243_1) );
	NOR2X1 NOR2X1_212 ( .A(_abc_3927_n892), .B(_abc_3927_n1243_1), .Y(_abc_3927_n1244) );
	NAND2X1 NAND2X1_343 ( .A(_abc_3927_n1244), .B(_abc_3927_n1242), .Y(_abc_3927_n1245_1) );
	XNOR2X1 XNOR2X1_42 ( .A(_abc_3927_n1206), .B(_abc_3927_n1001), .Y(_abc_3927_n1246) );
	NAND2X1 NAND2X1_344 ( .A(_abc_3927_n892), .B(_abc_3927_n1246), .Y(_abc_3927_n1247_1) );
	NAND2X1 NAND2X1_345 ( .A(_abc_3927_n1247_1), .B(_abc_3927_n1245_1), .Y(_abc_3927_n1248) );
	AND2X2 AND2X2_87 ( .A(_abc_3927_n1248), .B(_abc_3927_n365), .Y(currentaddr_20__FF_INPUT) );
	NOR2X1 NOR2X1_213 ( .A(_abc_3927_n1179), .B(_abc_3927_n815_1), .Y(_abc_3927_n1250) );
	NAND2X1 NAND2X1_346 ( .A(_abc_3927_n1180_1), .B(_abc_3927_n1250), .Y(_abc_3927_n1251_1) );
	NAND2X1 NAND2X1_347 ( .A(_abc_3927_n824), .B(_abc_3927_n1251_1), .Y(_abc_3927_n1252) );
	NAND2X1 NAND2X1_348 ( .A(_abc_3927_n1183), .B(_abc_3927_n1252), .Y(_abc_3927_n1253_1) );
	NAND2X1 NAND2X1_349 ( .A(_abc_3927_n405), .B(_abc_3927_n1253_1), .Y(_abc_3927_n1254) );
	NOR2X1 NOR2X1_214 ( .A(reg_fh_value_3_), .B(_abc_3927_n405), .Y(_abc_3927_n1255_1) );
	NOR2X1 NOR2X1_215 ( .A(_abc_3927_n892), .B(_abc_3927_n1255_1), .Y(_abc_3927_n1256) );
	NAND2X1 NAND2X1_350 ( .A(_abc_3927_n1256), .B(_abc_3927_n1254), .Y(_abc_3927_n1257_1) );
	NAND2X1 NAND2X1_351 ( .A(_abc_3927_n1024_1), .B(_abc_3927_n984), .Y(_abc_3927_n1258) );
	NAND2X1 NAND2X1_352 ( .A(_abc_3927_n1033), .B(_abc_3927_n1258), .Y(_abc_3927_n1259_1) );
	NAND2X1 NAND2X1_353 ( .A(_abc_3927_n1012), .B(_abc_3927_n1259_1), .Y(_abc_3927_n1260) );
	NAND2X1 NAND2X1_354 ( .A(_abc_3927_n1035), .B(_abc_3927_n1260), .Y(_abc_3927_n1261_1) );
	XOR2X1 XOR2X1_23 ( .A(_abc_3927_n1261_1), .B(_abc_3927_n1007), .Y(_abc_3927_n1262) );
	NAND2X1 NAND2X1_355 ( .A(_abc_3927_n892), .B(_abc_3927_n1262), .Y(_abc_3927_n1263_1) );
	NAND2X1 NAND2X1_356 ( .A(_abc_3927_n1263_1), .B(_abc_3927_n1257_1), .Y(_abc_3927_n1264) );
	AND2X2 AND2X2_88 ( .A(_abc_3927_n1264), .B(_abc_3927_n365), .Y(currentaddr_19__FF_INPUT) );
	NOR2X1 NOR2X1_216 ( .A(_abc_3927_n1008), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1266) );
	NAND2X1 NAND2X1_357 ( .A(_abc_3927_n825), .B(_abc_3927_n1106_1), .Y(_abc_3927_n1267_1) );
	XNOR2X1 XNOR2X1_43 ( .A(_abc_3927_n1267_1), .B(currentaddr_18_), .Y(_abc_3927_n1268) );
	AND2X2 AND2X2_89 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1268), .Y(_abc_3927_n1269_1) );
	NOR2X1 NOR2X1_217 ( .A(_abc_3927_n1266), .B(_abc_3927_n1269_1), .Y(_abc_3927_n1270) );
	NAND2X1 NAND2X1_358 ( .A(_abc_3927_n405), .B(_abc_3927_n1270), .Y(_abc_3927_n1271_1) );
	NOR2X1 NOR2X1_218 ( .A(reg_fh_value_2_), .B(_abc_3927_n405), .Y(_abc_3927_n1272) );
	NOR2X1 NOR2X1_219 ( .A(_abc_3927_n892), .B(_abc_3927_n1272), .Y(_abc_3927_n1273_1) );
	NAND2X1 NAND2X1_359 ( .A(_abc_3927_n1273_1), .B(_abc_3927_n1271_1), .Y(_abc_3927_n1274) );
	XOR2X1 XOR2X1_24 ( .A(_abc_3927_n1259_1), .B(_abc_3927_n1012), .Y(_abc_3927_n1275_1) );
	NAND2X1 NAND2X1_360 ( .A(_abc_3927_n892), .B(_abc_3927_n1275_1), .Y(_abc_3927_n1276) );
	NAND2X1 NAND2X1_361 ( .A(_abc_3927_n1276), .B(_abc_3927_n1274), .Y(_abc_3927_n1277_1) );
	AND2X2 AND2X2_90 ( .A(_abc_3927_n1277_1), .B(_abc_3927_n365), .Y(currentaddr_18__FF_INPUT) );
	NAND2X1 NAND2X1_362 ( .A(currentaddr_17_), .B(_abc_3927_n815_1), .Y(_abc_3927_n1279_1) );
	NAND2X1 NAND2X1_363 ( .A(currentaddr_16_), .B(_abc_3927_n1106_1), .Y(_abc_3927_n1280) );
	XNOR2X1 XNOR2X1_44 ( .A(_abc_3927_n1280), .B(currentaddr_17_), .Y(_abc_3927_n1281_1) );
	NAND2X1 NAND2X1_364 ( .A(_abc_3927_n1281_1), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1282) );
	AND2X2 AND2X2_91 ( .A(_abc_3927_n1279_1), .B(_abc_3927_n1282), .Y(_abc_3927_n1283_1) );
	NAND2X1 NAND2X1_365 ( .A(_abc_3927_n405), .B(_abc_3927_n1283_1), .Y(_abc_3927_n1284) );
	NOR2X1 NOR2X1_220 ( .A(reg_fh_value_1_), .B(_abc_3927_n405), .Y(_abc_3927_n1285) );
	NOR2X1 NOR2X1_221 ( .A(_abc_3927_n892), .B(_abc_3927_n1285), .Y(_abc_3927_n1286) );
	NAND2X1 NAND2X1_366 ( .A(_abc_3927_n1286), .B(_abc_3927_n1284), .Y(_abc_3927_n1287) );
	AND2X2 AND2X2_92 ( .A(_abc_3927_n984), .B(_abc_3927_n1018), .Y(_abc_3927_n1288) );
	NOR2X1 NOR2X1_222 ( .A(_abc_3927_n1016), .B(_abc_3927_n1288), .Y(_abc_3927_n1289) );
	XOR2X1 XOR2X1_25 ( .A(_abc_3927_n1289), .B(_abc_3927_n1023), .Y(_abc_3927_n1290) );
	NAND2X1 NAND2X1_367 ( .A(_abc_3927_n892), .B(_abc_3927_n1290), .Y(_abc_3927_n1291) );
	NAND2X1 NAND2X1_368 ( .A(_abc_3927_n1291), .B(_abc_3927_n1287), .Y(_abc_3927_n1292) );
	AND2X2 AND2X2_93 ( .A(_abc_3927_n1292), .B(_abc_3927_n365), .Y(currentaddr_17__FF_INPUT) );
	NAND2X1 NAND2X1_369 ( .A(_abc_3927_n831), .B(_abc_3927_n1250), .Y(_abc_3927_n1294) );
	XOR2X1 XOR2X1_26 ( .A(_abc_3927_n1294), .B(currentaddr_16_), .Y(_abc_3927_n1295) );
	NAND2X1 NAND2X1_370 ( .A(_abc_3927_n405), .B(_abc_3927_n1295), .Y(_abc_3927_n1296) );
	NOR2X1 NOR2X1_223 ( .A(reg_fh_value_0_), .B(_abc_3927_n405), .Y(_abc_3927_n1297) );
	NOR2X1 NOR2X1_224 ( .A(_abc_3927_n892), .B(_abc_3927_n1297), .Y(_abc_3927_n1298) );
	NAND2X1 NAND2X1_371 ( .A(_abc_3927_n1298), .B(_abc_3927_n1296), .Y(_abc_3927_n1299) );
	XNOR2X1 XNOR2X1_45 ( .A(_abc_3927_n984), .B(_abc_3927_n1019), .Y(_abc_3927_n1300) );
	NAND2X1 NAND2X1_372 ( .A(_abc_3927_n892), .B(_abc_3927_n1300), .Y(_abc_3927_n1301) );
	NAND2X1 NAND2X1_373 ( .A(_abc_3927_n1301), .B(_abc_3927_n1299), .Y(_abc_3927_n1302) );
	AND2X2 AND2X2_94 ( .A(_abc_3927_n1302), .B(_abc_3927_n365), .Y(currentaddr_16__FF_INPUT) );
	NAND2X1 NAND2X1_374 ( .A(currentaddr_14_), .B(_abc_3927_n1250), .Y(_abc_3927_n1304) );
	NAND2X1 NAND2X1_375 ( .A(_abc_3927_n829), .B(_abc_3927_n1304), .Y(_abc_3927_n1305) );
	NAND2X1 NAND2X1_376 ( .A(_abc_3927_n1294), .B(_abc_3927_n1305), .Y(_abc_3927_n1306) );
	NAND2X1 NAND2X1_377 ( .A(_abc_3927_n405), .B(_abc_3927_n1306), .Y(_abc_3927_n1307) );
	NOR2X1 NOR2X1_225 ( .A(reg_fl_value_15_), .B(_abc_3927_n405), .Y(_abc_3927_n1308) );
	NOR2X1 NOR2X1_226 ( .A(_abc_3927_n892), .B(_abc_3927_n1308), .Y(_abc_3927_n1309) );
	NAND2X1 NAND2X1_378 ( .A(_abc_3927_n1309), .B(_abc_3927_n1307), .Y(_abc_3927_n1310) );
	INVX1 INVX1_83 ( .A(_abc_3927_n950), .Y(_abc_3927_n1311) );
	INVX1 INVX1_84 ( .A(_abc_3927_n975_1), .Y(_abc_3927_n1312) );
	INVX1 INVX1_85 ( .A(_abc_3927_n965), .Y(_abc_3927_n1313) );
	NAND2X1 NAND2X1_379 ( .A(_abc_3927_n1313), .B(_abc_3927_n934_1), .Y(_abc_3927_n1314) );
	NAND2X1 NAND2X1_380 ( .A(_abc_3927_n1312), .B(_abc_3927_n1314), .Y(_abc_3927_n1315) );
	NAND2X1 NAND2X1_381 ( .A(_abc_3927_n1311), .B(_abc_3927_n1315), .Y(_abc_3927_n1316) );
	NAND2X1 NAND2X1_382 ( .A(_abc_3927_n978), .B(_abc_3927_n1316), .Y(_abc_3927_n1317) );
	AND2X2 AND2X2_95 ( .A(_abc_3927_n1317), .B(_abc_3927_n940_1), .Y(_abc_3927_n1318) );
	NOR2X1 NOR2X1_227 ( .A(_abc_3927_n938_1), .B(_abc_3927_n1318), .Y(_abc_3927_n1319) );
	XNOR2X1 XNOR2X1_46 ( .A(_abc_3927_n1319), .B(_abc_3927_n937_1), .Y(_abc_3927_n1320) );
	NAND2X1 NAND2X1_383 ( .A(_abc_3927_n892), .B(_abc_3927_n1320), .Y(_abc_3927_n1321) );
	NAND2X1 NAND2X1_384 ( .A(_abc_3927_n1321), .B(_abc_3927_n1310), .Y(_abc_3927_n1322) );
	AND2X2 AND2X2_96 ( .A(_abc_3927_n1322), .B(_abc_3927_n365), .Y(currentaddr_15__FF_INPUT) );
	XNOR2X1 XNOR2X1_47 ( .A(_abc_3927_n1250), .B(currentaddr_14_), .Y(_abc_3927_n1324) );
	NAND2X1 NAND2X1_385 ( .A(_abc_3927_n405), .B(_abc_3927_n1324), .Y(_abc_3927_n1325) );
	NOR2X1 NOR2X1_228 ( .A(reg_fl_value_14_), .B(_abc_3927_n405), .Y(_abc_3927_n1326) );
	NOR2X1 NOR2X1_229 ( .A(_abc_3927_n892), .B(_abc_3927_n1326), .Y(_abc_3927_n1327) );
	NAND2X1 NAND2X1_386 ( .A(_abc_3927_n1327), .B(_abc_3927_n1325), .Y(_abc_3927_n1328) );
	XOR2X1 XOR2X1_27 ( .A(_abc_3927_n1317), .B(_abc_3927_n940_1), .Y(_abc_3927_n1329) );
	NAND2X1 NAND2X1_387 ( .A(_abc_3927_n892), .B(_abc_3927_n1329), .Y(_abc_3927_n1330) );
	NAND2X1 NAND2X1_388 ( .A(_abc_3927_n1330), .B(_abc_3927_n1328), .Y(_abc_3927_n1331) );
	AND2X2 AND2X2_97 ( .A(_abc_3927_n1331), .B(_abc_3927_n365), .Y(currentaddr_14__FF_INPUT) );
	NOR2X1 NOR2X1_230 ( .A(_abc_3927_n832), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1333_1) );
	INVX1 INVX1_86 ( .A(_abc_3927_n1100_1), .Y(_abc_3927_n1334_1) );
	NOR2X1 NOR2X1_231 ( .A(_abc_3927_n1105), .B(_abc_3927_n1334_1), .Y(_abc_3927_n1335_1) );
	NAND2X1 NAND2X1_389 ( .A(currentaddr_12_), .B(_abc_3927_n1335_1), .Y(_abc_3927_n1336_1) );
	XNOR2X1 XNOR2X1_48 ( .A(_abc_3927_n1336_1), .B(currentaddr_13_), .Y(_abc_3927_n1337_1) );
	AND2X2 AND2X2_98 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1337_1), .Y(_abc_3927_n1338_1) );
	NOR2X1 NOR2X1_232 ( .A(_abc_3927_n1333_1), .B(_abc_3927_n1338_1), .Y(_abc_3927_n1339_1) );
	NAND2X1 NAND2X1_390 ( .A(_abc_3927_n405), .B(_abc_3927_n1339_1), .Y(_abc_3927_n1340_1) );
	NOR2X1 NOR2X1_233 ( .A(reg_fl_value_13_), .B(_abc_3927_n405), .Y(_abc_3927_n1341_1) );
	NOR2X1 NOR2X1_234 ( .A(_abc_3927_n892), .B(_abc_3927_n1341_1), .Y(_abc_3927_n1342_1) );
	NAND2X1 NAND2X1_391 ( .A(_abc_3927_n1342_1), .B(_abc_3927_n1340_1), .Y(_abc_3927_n1343_1) );
	NAND2X1 NAND2X1_392 ( .A(_abc_3927_n945_1), .B(_abc_3927_n1315), .Y(_abc_3927_n1344_1) );
	NAND2X1 NAND2X1_393 ( .A(_abc_3927_n942_1), .B(_abc_3927_n1344_1), .Y(_abc_3927_n1345_1) );
	XNOR2X1 XNOR2X1_49 ( .A(_abc_3927_n1345_1), .B(_abc_3927_n949), .Y(_abc_3927_n1346_1) );
	NAND2X1 NAND2X1_394 ( .A(_abc_3927_n892), .B(_abc_3927_n1346_1), .Y(_abc_3927_n1347_1) );
	NAND2X1 NAND2X1_395 ( .A(_abc_3927_n1347_1), .B(_abc_3927_n1343_1), .Y(_abc_3927_n1348) );
	AND2X2 AND2X2_99 ( .A(_abc_3927_n1348), .B(_abc_3927_n365), .Y(currentaddr_13__FF_INPUT) );
	NOR2X1 NOR2X1_235 ( .A(_abc_3927_n833), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1350) );
	XNOR2X1 XNOR2X1_50 ( .A(_abc_3927_n1335_1), .B(_abc_3927_n833), .Y(_abc_3927_n1351) );
	AND2X2 AND2X2_100 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1351), .Y(_abc_3927_n1352) );
	NOR2X1 NOR2X1_236 ( .A(_abc_3927_n1350), .B(_abc_3927_n1352), .Y(_abc_3927_n1353) );
	NAND2X1 NAND2X1_396 ( .A(_abc_3927_n405), .B(_abc_3927_n1353), .Y(_abc_3927_n1354) );
	NOR2X1 NOR2X1_237 ( .A(reg_fl_value_12_), .B(_abc_3927_n405), .Y(_abc_3927_n1355) );
	NOR2X1 NOR2X1_238 ( .A(_abc_3927_n892), .B(_abc_3927_n1355), .Y(_abc_3927_n1356) );
	NAND2X1 NAND2X1_397 ( .A(_abc_3927_n1356), .B(_abc_3927_n1354), .Y(_abc_3927_n1357) );
	XNOR2X1 XNOR2X1_51 ( .A(_abc_3927_n1315), .B(_abc_3927_n946_1), .Y(_abc_3927_n1358) );
	NAND2X1 NAND2X1_398 ( .A(_abc_3927_n892), .B(_abc_3927_n1358), .Y(_abc_3927_n1359) );
	NAND2X1 NAND2X1_399 ( .A(_abc_3927_n1359), .B(_abc_3927_n1357), .Y(_abc_3927_n1360) );
	AND2X2 AND2X2_101 ( .A(_abc_3927_n1360), .B(_abc_3927_n365), .Y(currentaddr_12__FF_INPUT) );
	NOR2X1 NOR2X1_239 ( .A(_abc_3927_n836), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1362) );
	NOR2X1 NOR2X1_240 ( .A(_abc_3927_n851), .B(_abc_3927_n1105), .Y(_abc_3927_n1363) );
	NAND2X1 NAND2X1_400 ( .A(currentaddr_10_), .B(_abc_3927_n1363), .Y(_abc_3927_n1364) );
	XNOR2X1 XNOR2X1_52 ( .A(_abc_3927_n1364), .B(currentaddr_11_), .Y(_abc_3927_n1365) );
	AND2X2 AND2X2_102 ( .A(_abc_3927_n1094_1), .B(_abc_3927_n1365), .Y(_abc_3927_n1366) );
	NOR2X1 NOR2X1_241 ( .A(_abc_3927_n1362), .B(_abc_3927_n1366), .Y(_abc_3927_n1367) );
	NAND2X1 NAND2X1_401 ( .A(_abc_3927_n405), .B(_abc_3927_n1367), .Y(_abc_3927_n1368) );
	NOR2X1 NOR2X1_242 ( .A(reg_fl_value_11_), .B(_abc_3927_n405), .Y(_abc_3927_n1369) );
	NOR2X1 NOR2X1_243 ( .A(_abc_3927_n892), .B(_abc_3927_n1369), .Y(_abc_3927_n1370) );
	NAND2X1 NAND2X1_402 ( .A(_abc_3927_n1370), .B(_abc_3927_n1368), .Y(_abc_3927_n1371) );
	NAND2X1 NAND2X1_403 ( .A(_abc_3927_n963), .B(_abc_3927_n934_1), .Y(_abc_3927_n1372) );
	NAND2X1 NAND2X1_404 ( .A(_abc_3927_n970), .B(_abc_3927_n1372), .Y(_abc_3927_n1373) );
	NAND2X1 NAND2X1_405 ( .A(_abc_3927_n955), .B(_abc_3927_n1373), .Y(_abc_3927_n1374) );
	NAND2X1 NAND2X1_406 ( .A(_abc_3927_n972_1), .B(_abc_3927_n1374), .Y(_abc_3927_n1375) );
	XOR2X1 XOR2X1_28 ( .A(_abc_3927_n1375), .B(_abc_3927_n954), .Y(_abc_3927_n1376) );
	NAND2X1 NAND2X1_407 ( .A(_abc_3927_n892), .B(_abc_3927_n1376), .Y(_abc_3927_n1377) );
	NAND2X1 NAND2X1_408 ( .A(_abc_3927_n1377), .B(_abc_3927_n1371), .Y(_abc_3927_n1378) );
	AND2X2 AND2X2_103 ( .A(_abc_3927_n1378), .B(_abc_3927_n365), .Y(currentaddr_11__FF_INPUT) );
	NOR2X1 NOR2X1_244 ( .A(_abc_3927_n847), .B(_abc_3927_n815_1), .Y(_abc_3927_n1380_1) );
	NAND2X1 NAND2X1_409 ( .A(_abc_3927_n850), .B(_abc_3927_n1380_1), .Y(_abc_3927_n1381_1) );
	XNOR2X1 XNOR2X1_53 ( .A(_abc_3927_n1381_1), .B(_abc_3927_n837), .Y(_abc_3927_n1382_1) );
	NAND2X1 NAND2X1_410 ( .A(_abc_3927_n405), .B(_abc_3927_n1382_1), .Y(_abc_3927_n1383_1) );
	NOR2X1 NOR2X1_245 ( .A(reg_fl_value_10_), .B(_abc_3927_n405), .Y(_abc_3927_n1384_1) );
	NOR2X1 NOR2X1_246 ( .A(_abc_3927_n892), .B(_abc_3927_n1384_1), .Y(_abc_3927_n1385_1) );
	NAND2X1 NAND2X1_411 ( .A(_abc_3927_n1385_1), .B(_abc_3927_n1383_1), .Y(_abc_3927_n1386_1) );
	XOR2X1 XOR2X1_29 ( .A(_abc_3927_n1373), .B(_abc_3927_n955), .Y(_abc_3927_n1387_1) );
	NAND2X1 NAND2X1_412 ( .A(_abc_3927_n892), .B(_abc_3927_n1387_1), .Y(_abc_3927_n1388_1) );
	NAND2X1 NAND2X1_413 ( .A(_abc_3927_n1388_1), .B(_abc_3927_n1386_1), .Y(_abc_3927_n1389_1) );
	AND2X2 AND2X2_104 ( .A(_abc_3927_n1389_1), .B(_abc_3927_n365), .Y(currentaddr_10__FF_INPUT) );
	NAND2X1 NAND2X1_414 ( .A(currentaddr_8_), .B(_abc_3927_n1380_1), .Y(_abc_3927_n1391_1) );
	XNOR2X1 XNOR2X1_54 ( .A(_abc_3927_n1391_1), .B(_abc_3927_n848), .Y(_abc_3927_n1392_1) );
	NAND2X1 NAND2X1_415 ( .A(_abc_3927_n405), .B(_abc_3927_n1392_1), .Y(_abc_3927_n1393_1) );
	NOR2X1 NOR2X1_247 ( .A(reg_fl_value_9_), .B(_abc_3927_n405), .Y(_abc_3927_n1394_1) );
	NOR2X1 NOR2X1_248 ( .A(_abc_3927_n892), .B(_abc_3927_n1394_1), .Y(_abc_3927_n1395) );
	NAND2X1 NAND2X1_416 ( .A(_abc_3927_n1395), .B(_abc_3927_n1393_1), .Y(_abc_3927_n1396) );
	INVX1 INVX1_87 ( .A(_abc_3927_n962), .Y(_abc_3927_n1397) );
	NAND2X1 NAND2X1_417 ( .A(_abc_3927_n1397), .B(_abc_3927_n934_1), .Y(_abc_3927_n1398) );
	NAND2X1 NAND2X1_418 ( .A(_abc_3927_n960), .B(_abc_3927_n1398), .Y(_abc_3927_n1399) );
	XNOR2X1 XNOR2X1_55 ( .A(_abc_3927_n1399), .B(_abc_3927_n959), .Y(_abc_3927_n1400) );
	NAND2X1 NAND2X1_419 ( .A(_abc_3927_n892), .B(_abc_3927_n1400), .Y(_abc_3927_n1401) );
	NAND2X1 NAND2X1_420 ( .A(_abc_3927_n1401), .B(_abc_3927_n1396), .Y(_abc_3927_n1402) );
	AND2X2 AND2X2_105 ( .A(_abc_3927_n1402), .B(_abc_3927_n365), .Y(currentaddr_9__FF_INPUT) );
	INVX1 INVX1_88 ( .A(_abc_3927_n1380_1), .Y(_abc_3927_n1404) );
	NAND2X1 NAND2X1_421 ( .A(_abc_3927_n849), .B(_abc_3927_n1404), .Y(_abc_3927_n1405) );
	NAND2X1 NAND2X1_422 ( .A(_abc_3927_n1391_1), .B(_abc_3927_n1405), .Y(_abc_3927_n1406) );
	NAND2X1 NAND2X1_423 ( .A(_abc_3927_n405), .B(_abc_3927_n1406), .Y(_abc_3927_n1407) );
	NOR2X1 NOR2X1_249 ( .A(reg_fl_value_8_), .B(_abc_3927_n405), .Y(_abc_3927_n1408) );
	NOR2X1 NOR2X1_250 ( .A(_abc_3927_n892), .B(_abc_3927_n1408), .Y(_abc_3927_n1409) );
	NAND2X1 NAND2X1_424 ( .A(_abc_3927_n1409), .B(_abc_3927_n1407), .Y(_abc_3927_n1410) );
	XNOR2X1 XNOR2X1_56 ( .A(_abc_3927_n934_1), .B(_abc_3927_n962), .Y(_abc_3927_n1411) );
	NAND2X1 NAND2X1_425 ( .A(_abc_3927_n892), .B(_abc_3927_n1411), .Y(_abc_3927_n1412) );
	NAND2X1 NAND2X1_426 ( .A(_abc_3927_n1412), .B(_abc_3927_n1410), .Y(_abc_3927_n1413) );
	AND2X2 AND2X2_106 ( .A(_abc_3927_n1413), .B(_abc_3927_n365), .Y(currentaddr_8__FF_INPUT) );
	NAND2X1 NAND2X1_427 ( .A(_abc_3927_n846), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1415) );
	XOR2X1 XOR2X1_30 ( .A(_abc_3927_n1415), .B(currentaddr_7_), .Y(_abc_3927_n1416) );
	NAND2X1 NAND2X1_428 ( .A(_abc_3927_n405), .B(_abc_3927_n1416), .Y(_abc_3927_n1417) );
	NOR2X1 NOR2X1_251 ( .A(reg_fl_value_7_), .B(_abc_3927_n405), .Y(_abc_3927_n1418) );
	NOR2X1 NOR2X1_252 ( .A(_abc_3927_n892), .B(_abc_3927_n1418), .Y(_abc_3927_n1419) );
	NAND2X1 NAND2X1_429 ( .A(_abc_3927_n1419), .B(_abc_3927_n1417), .Y(_abc_3927_n1420) );
	INVX1 INVX1_89 ( .A(_abc_3927_n916), .Y(_abc_3927_n1421) );
	INVX1 INVX1_90 ( .A(_abc_3927_n924), .Y(_abc_3927_n1422) );
	NAND2X1 NAND2X1_430 ( .A(_abc_3927_n1422), .B(_abc_3927_n912), .Y(_abc_3927_n1423) );
	NAND2X1 NAND2X1_431 ( .A(_abc_3927_n929), .B(_abc_3927_n1423), .Y(_abc_3927_n1424) );
	NAND2X1 NAND2X1_432 ( .A(_abc_3927_n918), .B(_abc_3927_n1424), .Y(_abc_3927_n1425_1) );
	NAND2X1 NAND2X1_433 ( .A(_abc_3927_n1421), .B(_abc_3927_n1425_1), .Y(_abc_3927_n1426_1) );
	XOR2X1 XOR2X1_31 ( .A(_abc_3927_n1426_1), .B(_abc_3927_n915), .Y(_abc_3927_n1427_1) );
	NAND2X1 NAND2X1_434 ( .A(_abc_3927_n892), .B(_abc_3927_n1427_1), .Y(_abc_3927_n1428_1) );
	NAND2X1 NAND2X1_435 ( .A(_abc_3927_n1428_1), .B(_abc_3927_n1420), .Y(_abc_3927_n1429_1) );
	AND2X2 AND2X2_107 ( .A(_abc_3927_n1429_1), .B(_abc_3927_n365), .Y(currentaddr_7__FF_INPUT) );
	NAND2X1 NAND2X1_436 ( .A(reg_fl_value_6_), .B(_abc_3927_n404), .Y(_abc_3927_n1431_1) );
	OR2X2 OR2X2_64 ( .A(_abc_3927_n815_1), .B(_abc_3927_n845), .Y(_abc_3927_n1432_1) );
	NAND2X1 NAND2X1_437 ( .A(_abc_3927_n839), .B(_abc_3927_n1432_1), .Y(_abc_3927_n1433_1) );
	AND2X2 AND2X2_108 ( .A(_abc_3927_n1433_1), .B(_abc_3927_n1415), .Y(_abc_3927_n1434_1) );
	NAND2X1 NAND2X1_438 ( .A(_abc_3927_n405), .B(_abc_3927_n1434_1), .Y(_abc_3927_n1435_1) );
	NAND2X1 NAND2X1_439 ( .A(_abc_3927_n1431_1), .B(_abc_3927_n1435_1), .Y(_abc_3927_n1436_1) );
	NOR2X1 NOR2X1_253 ( .A(_abc_3927_n892), .B(_abc_3927_n1436_1), .Y(_abc_3927_n1437_1) );
	XNOR2X1 XNOR2X1_57 ( .A(_abc_3927_n1424), .B(_abc_3927_n918), .Y(_abc_3927_n1438_1) );
	NAND2X1 NAND2X1_440 ( .A(_abc_3927_n892), .B(_abc_3927_n1438_1), .Y(_abc_3927_n1439_1) );
	NAND2X1 NAND2X1_441 ( .A(_abc_3927_n365), .B(_abc_3927_n1439_1), .Y(_abc_3927_n1440_1) );
	NOR2X1 NOR2X1_254 ( .A(_abc_3927_n1440_1), .B(_abc_3927_n1437_1), .Y(currentaddr_6__FF_INPUT) );
	NAND2X1 NAND2X1_442 ( .A(_abc_3927_n844), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1442) );
	XOR2X1 XOR2X1_32 ( .A(_abc_3927_n1442), .B(currentaddr_5_), .Y(_abc_3927_n1443) );
	NAND2X1 NAND2X1_443 ( .A(_abc_3927_n405), .B(_abc_3927_n1443), .Y(_abc_3927_n1444) );
	NOR2X1 NOR2X1_255 ( .A(reg_fl_value_5_), .B(_abc_3927_n405), .Y(_abc_3927_n1445) );
	NOR2X1 NOR2X1_256 ( .A(_abc_3927_n892), .B(_abc_3927_n1445), .Y(_abc_3927_n1446) );
	NAND2X1 NAND2X1_444 ( .A(_abc_3927_n1446), .B(_abc_3927_n1444), .Y(_abc_3927_n1447) );
	NAND2X1 NAND2X1_445 ( .A(_abc_3927_n920), .B(_abc_3927_n912), .Y(_abc_3927_n1448) );
	NAND2X1 NAND2X1_446 ( .A(_abc_3927_n927), .B(_abc_3927_n1448), .Y(_abc_3927_n1449) );
	XOR2X1 XOR2X1_33 ( .A(_abc_3927_n1449), .B(_abc_3927_n923), .Y(_abc_3927_n1450) );
	NAND2X1 NAND2X1_447 ( .A(_abc_3927_n892), .B(_abc_3927_n1450), .Y(_abc_3927_n1451) );
	NAND2X1 NAND2X1_448 ( .A(_abc_3927_n1451), .B(_abc_3927_n1447), .Y(_abc_3927_n1452) );
	AND2X2 AND2X2_109 ( .A(_abc_3927_n1452), .B(_abc_3927_n365), .Y(currentaddr_5__FF_INPUT) );
	NAND2X1 NAND2X1_449 ( .A(_abc_3927_n843), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1454) );
	XOR2X1 XOR2X1_34 ( .A(_abc_3927_n1454), .B(currentaddr_4_), .Y(_abc_3927_n1455) );
	NAND2X1 NAND2X1_450 ( .A(_abc_3927_n405), .B(_abc_3927_n1455), .Y(_abc_3927_n1456) );
	NOR2X1 NOR2X1_257 ( .A(reg_fl_value_4_), .B(_abc_3927_n405), .Y(_abc_3927_n1457) );
	NOR2X1 NOR2X1_258 ( .A(_abc_3927_n892), .B(_abc_3927_n1457), .Y(_abc_3927_n1458) );
	NAND2X1 NAND2X1_451 ( .A(_abc_3927_n1458), .B(_abc_3927_n1456), .Y(_abc_3927_n1459) );
	XOR2X1 XOR2X1_35 ( .A(_abc_3927_n912), .B(_abc_3927_n920), .Y(_abc_3927_n1460) );
	NAND2X1 NAND2X1_452 ( .A(_abc_3927_n892), .B(_abc_3927_n1460), .Y(_abc_3927_n1461) );
	NAND2X1 NAND2X1_453 ( .A(_abc_3927_n1461), .B(_abc_3927_n1459), .Y(_abc_3927_n1462) );
	AND2X2 AND2X2_110 ( .A(_abc_3927_n1462), .B(_abc_3927_n365), .Y(currentaddr_4__FF_INPUT) );
	NAND2X1 NAND2X1_454 ( .A(_abc_3927_n842), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1464) );
	XOR2X1 XOR2X1_36 ( .A(_abc_3927_n1464), .B(currentaddr_3_), .Y(_abc_3927_n1465) );
	NAND2X1 NAND2X1_455 ( .A(_abc_3927_n405), .B(_abc_3927_n1465), .Y(_abc_3927_n1466) );
	NOR2X1 NOR2X1_259 ( .A(reg_fl_value_3_), .B(_abc_3927_n405), .Y(_abc_3927_n1467) );
	NOR2X1 NOR2X1_260 ( .A(_abc_3927_n892), .B(_abc_3927_n1467), .Y(_abc_3927_n1468) );
	NAND2X1 NAND2X1_456 ( .A(_abc_3927_n1468), .B(_abc_3927_n1466), .Y(_abc_3927_n1469) );
	INVX1 INVX1_91 ( .A(_abc_3927_n902), .Y(_abc_3927_n1470) );
	NOR2X1 NOR2X1_261 ( .A(_abc_3927_n906), .B(_abc_3927_n1470), .Y(_abc_3927_n1471) );
	INVX1 INVX1_92 ( .A(_abc_3927_n1471), .Y(_abc_3927_n1472) );
	NAND2X1 NAND2X1_457 ( .A(_abc_3927_n904), .B(_abc_3927_n1472), .Y(_abc_3927_n1473) );
	XNOR2X1 XNOR2X1_58 ( .A(_abc_3927_n1473), .B(_abc_3927_n903), .Y(_abc_3927_n1474) );
	NAND2X1 NAND2X1_458 ( .A(_abc_3927_n892), .B(_abc_3927_n1474), .Y(_abc_3927_n1475) );
	NAND2X1 NAND2X1_459 ( .A(_abc_3927_n1475), .B(_abc_3927_n1469), .Y(_abc_3927_n1476) );
	AND2X2 AND2X2_111 ( .A(_abc_3927_n1476), .B(_abc_3927_n365), .Y(currentaddr_3__FF_INPUT) );
	NOR2X1 NOR2X1_262 ( .A(_abc_3927_n841), .B(_abc_3927_n815_1), .Y(_abc_3927_n1478) );
	XNOR2X1 XNOR2X1_59 ( .A(_abc_3927_n1478), .B(currentaddr_2_), .Y(_abc_3927_n1479_1) );
	NAND2X1 NAND2X1_460 ( .A(_abc_3927_n405), .B(_abc_3927_n1479_1), .Y(_abc_3927_n1480_1) );
	NOR2X1 NOR2X1_263 ( .A(reg_fl_value_2_), .B(_abc_3927_n405), .Y(_abc_3927_n1481_1) );
	NOR2X1 NOR2X1_264 ( .A(_abc_3927_n892), .B(_abc_3927_n1481_1), .Y(_abc_3927_n1482_1) );
	NAND2X1 NAND2X1_461 ( .A(_abc_3927_n1482_1), .B(_abc_3927_n1480_1), .Y(_abc_3927_n1483_1) );
	NAND2X1 NAND2X1_462 ( .A(_abc_3927_n906), .B(_abc_3927_n1470), .Y(_abc_3927_n1484_1) );
	NOR2X1 NOR2X1_265 ( .A(_abc_3927_n1471), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1485_1) );
	NAND2X1 NAND2X1_463 ( .A(_abc_3927_n1484_1), .B(_abc_3927_n1485_1), .Y(_abc_3927_n1486_1) );
	NAND2X1 NAND2X1_464 ( .A(_abc_3927_n1486_1), .B(_abc_3927_n1483_1), .Y(_abc_3927_n1487_1) );
	AND2X2 AND2X2_112 ( .A(_abc_3927_n1487_1), .B(_abc_3927_n365), .Y(currentaddr_2__FF_INPUT) );
	INVX1 INVX1_93 ( .A(currentaddr_1_), .Y(_abc_3927_n1489_1) );
	NAND2X1 NAND2X1_465 ( .A(currentaddr_0_), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1490_1) );
	NAND2X1 NAND2X1_466 ( .A(_abc_3927_n1489_1), .B(_abc_3927_n1490_1), .Y(_abc_3927_n1491_1) );
	NOR2X1 NOR2X1_266 ( .A(_abc_3927_n404), .B(_abc_3927_n1478), .Y(_abc_3927_n1492_1) );
	NAND2X1 NAND2X1_467 ( .A(_abc_3927_n1491_1), .B(_abc_3927_n1492_1), .Y(_abc_3927_n1493_1) );
	NAND2X1 NAND2X1_468 ( .A(reg_fl_value_1_), .B(_abc_3927_n404), .Y(_abc_3927_n1494_1) );
	NAND2X1 NAND2X1_469 ( .A(_abc_3927_n1494_1), .B(_abc_3927_n1493_1), .Y(_abc_3927_n1495) );
	NOR2X1 NOR2X1_267 ( .A(_abc_3927_n892), .B(_abc_3927_n1495), .Y(_abc_3927_n1496) );
	XNOR2X1 XNOR2X1_60 ( .A(_abc_3927_n900), .B(_abc_3927_n898), .Y(_abc_3927_n1497) );
	NAND2X1 NAND2X1_470 ( .A(_abc_3927_n1497), .B(_abc_3927_n892), .Y(_abc_3927_n1498) );
	NAND2X1 NAND2X1_471 ( .A(_abc_3927_n365), .B(_abc_3927_n1498), .Y(_abc_3927_n1499) );
	NOR2X1 NOR2X1_268 ( .A(_abc_3927_n1499), .B(_abc_3927_n1496), .Y(currentaddr_1__FF_INPUT) );
	NOR2X1 NOR2X1_269 ( .A(currentaddr_0_), .B(reg_sl_value_0_), .Y(_abc_3927_n1501) );
	NOR2X1 NOR2X1_270 ( .A(_abc_3927_n1501), .B(_abc_3927_n898), .Y(_abc_3927_n1502) );
	NAND2X1 NAND2X1_472 ( .A(_abc_3927_n1502), .B(_abc_3927_n892), .Y(_abc_3927_n1503) );
	XNOR2X1 XNOR2X1_61 ( .A(_abc_3927_n1094_1), .B(currentaddr_0_), .Y(_abc_3927_n1504_1) );
	NAND2X1 NAND2X1_473 ( .A(_abc_3927_n405), .B(_abc_3927_n1504_1), .Y(_abc_3927_n1505) );
	NOR2X1 NOR2X1_271 ( .A(reg_fl_value_0_), .B(_abc_3927_n405), .Y(_abc_3927_n1506_1) );
	NOR2X1 NOR2X1_272 ( .A(_abc_3927_n892), .B(_abc_3927_n1506_1), .Y(_abc_3927_n1507) );
	NAND2X1 NAND2X1_474 ( .A(_abc_3927_n1507), .B(_abc_3927_n1505), .Y(_abc_3927_n1508_1) );
	NAND2X1 NAND2X1_475 ( .A(_abc_3927_n1503), .B(_abc_3927_n1508_1), .Y(_abc_3927_n1509) );
	AND2X2 AND2X2_113 ( .A(_abc_3927_n1509), .B(_abc_3927_n365), .Y(currentaddr_0__FF_INPUT) );
	NAND2X1 NAND2X1_476 ( .A(_abc_3927_n365), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1511) );
	NOR2X1 NOR2X1_273 ( .A(_abc_3927_n583), .B(_abc_3927_n585), .Y(_abc_3927_n1512_1) );
	INVX1 INVX1_94 ( .A(_abc_3927_n1512_1), .Y(_abc_3927_n1513) );
	NOR2X1 NOR2X1_274 ( .A(_abc_3927_n591), .B(_abc_3927_n1513), .Y(_abc_3927_n1514) );
	NAND2X1 NAND2X1_477 ( .A(currentcol_3_), .B(_abc_3927_n1514), .Y(_abc_3927_n1515) );
	NOR2X1 NOR2X1_275 ( .A(_abc_3927_n569), .B(_abc_3927_n1515), .Y(_abc_3927_n1516) );
	NAND2X1 NAND2X1_478 ( .A(currentcol_5_), .B(_abc_3927_n1516), .Y(_abc_3927_n1517) );
	NOR2X1 NOR2X1_276 ( .A(_abc_3927_n562), .B(_abc_3927_n1517), .Y(_abc_3927_n1518_1) );
	NAND2X1 NAND2X1_479 ( .A(currentcol_7_), .B(_abc_3927_n1518_1), .Y(_abc_3927_n1519) );
	NOR2X1 NOR2X1_277 ( .A(_abc_3927_n548), .B(_abc_3927_n1519), .Y(_abc_3927_n1520) );
	NAND2X1 NAND2X1_480 ( .A(currentcol_9_), .B(_abc_3927_n1520), .Y(_abc_3927_n1521_1) );
	NOR2X1 NOR2X1_278 ( .A(_abc_3927_n604), .B(_abc_3927_n1521_1), .Y(_abc_3927_n1522_1) );
	NAND2X1 NAND2X1_481 ( .A(currentcol_11_), .B(_abc_3927_n1522_1), .Y(_abc_3927_n1523_1) );
	NOR2X1 NOR2X1_279 ( .A(_abc_3927_n531), .B(_abc_3927_n1523_1), .Y(_abc_3927_n1524) );
	NAND2X1 NAND2X1_482 ( .A(currentcol_13_), .B(_abc_3927_n1524), .Y(_abc_3927_n1525_1) );
	XNOR2X1 XNOR2X1_62 ( .A(_abc_3927_n1525_1), .B(_abc_3927_n524), .Y(_abc_3927_n1526) );
	NOR2X1 NOR2X1_280 ( .A(_abc_3927_n1511), .B(_abc_3927_n1526), .Y(currentcol_14__FF_INPUT) );
	INVX1 INVX1_95 ( .A(_abc_3927_n1524), .Y(_abc_3927_n1528_1) );
	NAND2X1 NAND2X1_483 ( .A(_abc_3927_n529), .B(_abc_3927_n1528_1), .Y(_abc_3927_n1529) );
	NAND2X1 NAND2X1_484 ( .A(_abc_3927_n1525_1), .B(_abc_3927_n1529), .Y(_abc_3927_n1530_1) );
	NOR2X1 NOR2X1_281 ( .A(_abc_3927_n1511), .B(_abc_3927_n1530_1), .Y(currentcol_13__FF_INPUT) );
	NAND2X1 NAND2X1_485 ( .A(_abc_3927_n531), .B(_abc_3927_n1523_1), .Y(_abc_3927_n1532) );
	NAND2X1 NAND2X1_486 ( .A(_abc_3927_n1532), .B(_abc_3927_n1528_1), .Y(_abc_3927_n1533) );
	NOR2X1 NOR2X1_282 ( .A(_abc_3927_n1511), .B(_abc_3927_n1533), .Y(currentcol_12__FF_INPUT) );
	INVX1 INVX1_96 ( .A(_abc_3927_n1522_1), .Y(_abc_3927_n1535) );
	NAND2X1 NAND2X1_487 ( .A(_abc_3927_n539), .B(_abc_3927_n1535), .Y(_abc_3927_n1536) );
	NAND2X1 NAND2X1_488 ( .A(_abc_3927_n1523_1), .B(_abc_3927_n1536), .Y(_abc_3927_n1537) );
	NOR2X1 NOR2X1_283 ( .A(_abc_3927_n1511), .B(_abc_3927_n1537), .Y(currentcol_11__FF_INPUT) );
	NAND2X1 NAND2X1_489 ( .A(_abc_3927_n604), .B(_abc_3927_n1521_1), .Y(_abc_3927_n1539) );
	NAND2X1 NAND2X1_490 ( .A(_abc_3927_n1539), .B(_abc_3927_n1535), .Y(_abc_3927_n1540) );
	NOR2X1 NOR2X1_284 ( .A(_abc_3927_n1511), .B(_abc_3927_n1540), .Y(currentcol_10__FF_INPUT) );
	INVX1 INVX1_97 ( .A(_abc_3927_n1520), .Y(_abc_3927_n1542) );
	NAND2X1 NAND2X1_491 ( .A(_abc_3927_n546), .B(_abc_3927_n1542), .Y(_abc_3927_n1543) );
	NAND2X1 NAND2X1_492 ( .A(_abc_3927_n1521_1), .B(_abc_3927_n1543), .Y(_abc_3927_n1544) );
	NOR2X1 NOR2X1_285 ( .A(_abc_3927_n1511), .B(_abc_3927_n1544), .Y(currentcol_9__FF_INPUT) );
	NAND2X1 NAND2X1_493 ( .A(_abc_3927_n548), .B(_abc_3927_n1519), .Y(_abc_3927_n1546) );
	NAND2X1 NAND2X1_494 ( .A(_abc_3927_n1546), .B(_abc_3927_n1542), .Y(_abc_3927_n1547) );
	NOR2X1 NOR2X1_286 ( .A(_abc_3927_n1511), .B(_abc_3927_n1547), .Y(currentcol_8__FF_INPUT) );
	INVX1 INVX1_98 ( .A(_abc_3927_n1518_1), .Y(_abc_3927_n1549) );
	NAND2X1 NAND2X1_495 ( .A(_abc_3927_n663), .B(_abc_3927_n1549), .Y(_abc_3927_n1550) );
	NAND2X1 NAND2X1_496 ( .A(_abc_3927_n1519), .B(_abc_3927_n1550), .Y(_abc_3927_n1551) );
	NOR2X1 NOR2X1_287 ( .A(_abc_3927_n1511), .B(_abc_3927_n1551), .Y(currentcol_7__FF_INPUT) );
	NAND2X1 NAND2X1_497 ( .A(_abc_3927_n562), .B(_abc_3927_n1517), .Y(_abc_3927_n1553) );
	NAND2X1 NAND2X1_498 ( .A(_abc_3927_n1553), .B(_abc_3927_n1549), .Y(_abc_3927_n1554) );
	NOR2X1 NOR2X1_288 ( .A(_abc_3927_n1511), .B(_abc_3927_n1554), .Y(currentcol_6__FF_INPUT) );
	INVX1 INVX1_99 ( .A(_abc_3927_n1516), .Y(_abc_3927_n1556) );
	NAND2X1 NAND2X1_499 ( .A(_abc_3927_n567), .B(_abc_3927_n1556), .Y(_abc_3927_n1557) );
	NAND2X1 NAND2X1_500 ( .A(_abc_3927_n1517), .B(_abc_3927_n1557), .Y(_abc_3927_n1558) );
	NOR2X1 NOR2X1_289 ( .A(_abc_3927_n1558), .B(_abc_3927_n1511), .Y(currentcol_5__FF_INPUT) );
	NAND2X1 NAND2X1_501 ( .A(_abc_3927_n569), .B(_abc_3927_n1515), .Y(_abc_3927_n1560) );
	NAND2X1 NAND2X1_502 ( .A(_abc_3927_n1560), .B(_abc_3927_n1556), .Y(_abc_3927_n1561) );
	NOR2X1 NOR2X1_290 ( .A(_abc_3927_n1561), .B(_abc_3927_n1511), .Y(currentcol_4__FF_INPUT) );
	XNOR2X1 XNOR2X1_63 ( .A(_abc_3927_n1514), .B(currentcol_3_), .Y(_abc_3927_n1563) );
	NOR2X1 NOR2X1_291 ( .A(_abc_3927_n1563), .B(_abc_3927_n1511), .Y(currentcol_3__FF_INPUT) );
	XNOR2X1 XNOR2X1_64 ( .A(_abc_3927_n1512_1), .B(currentcol_2_), .Y(_abc_3927_n1565) );
	NOR2X1 NOR2X1_292 ( .A(_abc_3927_n1565), .B(_abc_3927_n1511), .Y(currentcol_2__FF_INPUT) );
	NAND2X1 NAND2X1_503 ( .A(_abc_3927_n583), .B(_abc_3927_n585), .Y(_abc_3927_n1567) );
	NAND2X1 NAND2X1_504 ( .A(_abc_3927_n1567), .B(_abc_3927_n1513), .Y(_abc_3927_n1568) );
	NOR2X1 NOR2X1_293 ( .A(_abc_3927_n1568), .B(_abc_3927_n1511), .Y(currentcol_1__FF_INPUT) );
	NOR2X1 NOR2X1_294 ( .A(currentcol_0_), .B(_abc_3927_n1511), .Y(currentcol_0__FF_INPUT) );
	NOR2X1 NOR2X1_295 ( .A(reset), .B(_abc_3927_n404), .Y(_abc_3927_n1571) );
	INVX4 INVX4_3 ( .A(_abc_3927_n1571), .Y(_abc_3927_n1572) );
	NAND2X1 NAND2X1_505 ( .A(currentrow_0_), .B(currentrow_1_), .Y(_abc_3927_n1573) );
	NOR2X1 NOR2X1_296 ( .A(_abc_3927_n486_1), .B(_abc_3927_n1573), .Y(_abc_3927_n1574) );
	NAND2X1 NAND2X1_506 ( .A(currentrow_3_), .B(_abc_3927_n1574), .Y(_abc_3927_n1575) );
	NOR2X1 NOR2X1_297 ( .A(_abc_3927_n464), .B(_abc_3927_n1575), .Y(_abc_3927_n1576) );
	NAND2X1 NAND2X1_507 ( .A(currentrow_5_), .B(_abc_3927_n1576), .Y(_abc_3927_n1577) );
	NOR2X1 NOR2X1_298 ( .A(_abc_3927_n496), .B(_abc_3927_n1577), .Y(_abc_3927_n1578) );
	NAND2X1 NAND2X1_508 ( .A(currentrow_7_), .B(_abc_3927_n1578), .Y(_abc_3927_n1579) );
	NOR2X1 NOR2X1_299 ( .A(_abc_3927_n742), .B(_abc_3927_n1579), .Y(_abc_3927_n1580) );
	NAND2X1 NAND2X1_509 ( .A(currentrow_9_), .B(_abc_3927_n1580), .Y(_abc_3927_n1581) );
	NOR2X1 NOR2X1_300 ( .A(_abc_3927_n506), .B(_abc_3927_n1581), .Y(_abc_3927_n1582) );
	NAND2X1 NAND2X1_510 ( .A(currentrow_11_), .B(_abc_3927_n1582), .Y(_abc_3927_n1583) );
	NOR2X1 NOR2X1_301 ( .A(_abc_3927_n428_1), .B(_abc_3927_n1583), .Y(_abc_3927_n1584) );
	NAND2X1 NAND2X1_511 ( .A(currentrow_13_), .B(_abc_3927_n1584), .Y(_abc_3927_n1585) );
	NOR2X1 NOR2X1_302 ( .A(_abc_3927_n1088_1), .B(_abc_3927_n1585), .Y(_abc_3927_n1586) );
	XNOR2X1 XNOR2X1_65 ( .A(_abc_3927_n1586), .B(currentrow_14_), .Y(_abc_3927_n1587) );
	NOR2X1 NOR2X1_303 ( .A(_abc_3927_n1572), .B(_abc_3927_n1587), .Y(currentrow_14__FF_INPUT) );
	NAND2X1 NAND2X1_512 ( .A(_abc_3927_n892), .B(_abc_3927_n1584), .Y(_abc_3927_n1589) );
	XNOR2X1 XNOR2X1_66 ( .A(_abc_3927_n1589), .B(_abc_3927_n432_1), .Y(_abc_3927_n1590) );
	NOR2X1 NOR2X1_304 ( .A(_abc_3927_n1572), .B(_abc_3927_n1590), .Y(currentrow_13__FF_INPUT) );
	NOR2X1 NOR2X1_305 ( .A(_abc_3927_n1088_1), .B(_abc_3927_n1583), .Y(_abc_3927_n1592) );
	XNOR2X1 XNOR2X1_67 ( .A(_abc_3927_n1592), .B(currentrow_12_), .Y(_abc_3927_n1593) );
	NOR2X1 NOR2X1_306 ( .A(_abc_3927_n1572), .B(_abc_3927_n1593), .Y(currentrow_12__FF_INPUT) );
	NAND2X1 NAND2X1_513 ( .A(_abc_3927_n892), .B(_abc_3927_n1582), .Y(_abc_3927_n1595) );
	XNOR2X1 XNOR2X1_68 ( .A(_abc_3927_n1595), .B(_abc_3927_n438_1), .Y(_abc_3927_n1596) );
	NOR2X1 NOR2X1_307 ( .A(_abc_3927_n1572), .B(_abc_3927_n1596), .Y(currentrow_11__FF_INPUT) );
	NOR2X1 NOR2X1_308 ( .A(_abc_3927_n1088_1), .B(_abc_3927_n1581), .Y(_abc_3927_n1598) );
	XNOR2X1 XNOR2X1_69 ( .A(_abc_3927_n1598), .B(currentrow_10_), .Y(_abc_3927_n1599) );
	NOR2X1 NOR2X1_309 ( .A(_abc_3927_n1572), .B(_abc_3927_n1599), .Y(currentrow_10__FF_INPUT) );
	NAND2X1 NAND2X1_514 ( .A(_abc_3927_n892), .B(_abc_3927_n1580), .Y(_abc_3927_n1601) );
	XNOR2X1 XNOR2X1_70 ( .A(_abc_3927_n1601), .B(_abc_3927_n446), .Y(_abc_3927_n1602) );
	NOR2X1 NOR2X1_310 ( .A(_abc_3927_n1602), .B(_abc_3927_n1572), .Y(currentrow_9__FF_INPUT) );
	NOR2X1 NOR2X1_311 ( .A(_abc_3927_n1579), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1604) );
	XNOR2X1 XNOR2X1_71 ( .A(_abc_3927_n1604), .B(currentrow_8_), .Y(_abc_3927_n1605) );
	NOR2X1 NOR2X1_312 ( .A(_abc_3927_n1605), .B(_abc_3927_n1572), .Y(currentrow_8__FF_INPUT) );
	NAND2X1 NAND2X1_515 ( .A(_abc_3927_n1578), .B(_abc_3927_n892), .Y(_abc_3927_n1607) );
	XNOR2X1 XNOR2X1_72 ( .A(_abc_3927_n1607), .B(_abc_3927_n456), .Y(_abc_3927_n1608) );
	NOR2X1 NOR2X1_313 ( .A(_abc_3927_n1608), .B(_abc_3927_n1572), .Y(currentrow_7__FF_INPUT) );
	NOR2X1 NOR2X1_314 ( .A(_abc_3927_n1577), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1610) );
	XNOR2X1 XNOR2X1_73 ( .A(_abc_3927_n1610), .B(currentrow_6_), .Y(_abc_3927_n1611) );
	NOR2X1 NOR2X1_315 ( .A(_abc_3927_n1611), .B(_abc_3927_n1572), .Y(currentrow_6__FF_INPUT) );
	NAND2X1 NAND2X1_516 ( .A(_abc_3927_n1576), .B(_abc_3927_n892), .Y(_abc_3927_n1613) );
	XNOR2X1 XNOR2X1_74 ( .A(_abc_3927_n1613), .B(_abc_3927_n462), .Y(_abc_3927_n1614) );
	NOR2X1 NOR2X1_316 ( .A(_abc_3927_n1614), .B(_abc_3927_n1572), .Y(currentrow_5__FF_INPUT) );
	NOR2X1 NOR2X1_317 ( .A(_abc_3927_n1575), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1616) );
	XNOR2X1 XNOR2X1_75 ( .A(_abc_3927_n1616), .B(currentrow_4_), .Y(_abc_3927_n1617) );
	NOR2X1 NOR2X1_318 ( .A(_abc_3927_n1617), .B(_abc_3927_n1572), .Y(currentrow_4__FF_INPUT) );
	NAND2X1 NAND2X1_517 ( .A(_abc_3927_n1574), .B(_abc_3927_n892), .Y(_abc_3927_n1619) );
	XNOR2X1 XNOR2X1_76 ( .A(_abc_3927_n1619), .B(_abc_3927_n472), .Y(_abc_3927_n1620) );
	NOR2X1 NOR2X1_319 ( .A(_abc_3927_n1620), .B(_abc_3927_n1572), .Y(currentrow_3__FF_INPUT) );
	OR2X2 OR2X2_65 ( .A(_abc_3927_n1088_1), .B(_abc_3927_n1573), .Y(_abc_3927_n1622) );
	XNOR2X1 XNOR2X1_77 ( .A(_abc_3927_n1622), .B(_abc_3927_n486_1), .Y(_abc_3927_n1623) );
	NOR2X1 NOR2X1_320 ( .A(_abc_3927_n1623), .B(_abc_3927_n1572), .Y(currentrow_2__FF_INPUT) );
	NOR2X1 NOR2X1_321 ( .A(_abc_3927_n480_1), .B(_abc_3927_n1088_1), .Y(_abc_3927_n1625) );
	NOR2X1 NOR2X1_322 ( .A(currentrow_1_), .B(_abc_3927_n1625), .Y(_abc_3927_n1626) );
	NAND2X1 NAND2X1_518 ( .A(_abc_3927_n1622), .B(_abc_3927_n1571), .Y(_abc_3927_n1627) );
	NOR2X1 NOR2X1_323 ( .A(_abc_3927_n1626), .B(_abc_3927_n1627), .Y(currentrow_1__FF_INPUT) );
	NOR2X1 NOR2X1_324 ( .A(currentrow_0_), .B(_abc_3927_n892), .Y(_abc_3927_n1629) );
	NOR2X1 NOR2X1_325 ( .A(_abc_3927_n1629), .B(_abc_3927_n1625), .Y(_abc_3927_n1630) );
	AND2X2 AND2X2_114 ( .A(_abc_3927_n1571), .B(_abc_3927_n1630), .Y(currentrow_0__FF_INPUT) );
	NAND2X1 NAND2X1_519 ( .A(currentaddr_31_), .B(_abc_3927_n815_1), .Y(_abc_3927_n1632) );
	NAND2X1 NAND2X1_520 ( .A(_abc_3927_n409), .B(_abc_3927_n1108_1), .Y(_abc_3927_n1633) );
	NOR2X1 NOR2X1_326 ( .A(_abc_3927_n406), .B(_abc_3927_n1633), .Y(_abc_3927_n1634) );
	XOR2X1 XOR2X1_37 ( .A(_abc_3927_n1634), .B(currentaddr_31_), .Y(_abc_3927_n1635) );
	NAND2X1 NAND2X1_521 ( .A(_abc_3927_n1635), .B(_abc_3927_n1094_1), .Y(_abc_3927_n1636) );
	AND2X2 AND2X2_115 ( .A(_abc_3927_n1632), .B(_abc_3927_n1636), .Y(_abc_3927_n1637) );
	NAND2X1 NAND2X1_522 ( .A(_abc_3927_n405), .B(_abc_3927_n1637), .Y(_abc_3927_n1638) );
	NOR2X1 NOR2X1_327 ( .A(reg_fh_value_15_), .B(_abc_3927_n405), .Y(_abc_3927_n1639) );
	NOR2X1 NOR2X1_328 ( .A(_abc_3927_n892), .B(_abc_3927_n1639), .Y(_abc_3927_n1640) );
	NAND2X1 NAND2X1_523 ( .A(_abc_3927_n1640), .B(_abc_3927_n1638), .Y(_abc_3927_n1641) );
	NAND2X1 NAND2X1_524 ( .A(currentaddr_30_), .B(reg_sh_value_14_), .Y(_abc_3927_n1642) );
	NAND2X1 NAND2X1_525 ( .A(_abc_3927_n1642), .B(_abc_3927_n1087), .Y(_abc_3927_n1643) );
	XNOR2X1 XNOR2X1_78 ( .A(currentaddr_31_), .B(reg_sh_value_15_), .Y(_abc_3927_n1644) );
	XNOR2X1 XNOR2X1_79 ( .A(_abc_3927_n1643), .B(_abc_3927_n1644), .Y(_abc_3927_n1645) );
	NAND2X1 NAND2X1_526 ( .A(_abc_3927_n892), .B(_abc_3927_n1645), .Y(_abc_3927_n1646) );
	NAND2X1 NAND2X1_527 ( .A(_abc_3927_n1641), .B(_abc_3927_n1646), .Y(_abc_3927_n1647) );
	AND2X2 AND2X2_116 ( .A(_abc_3927_n1647), .B(_abc_3927_n365), .Y(currentaddr_31__FF_INPUT) );
	NOR2X1 NOR2X1_329 ( .A(_abc_3927_n524), .B(_abc_3927_n1525_1), .Y(_abc_3927_n1649) );
	XNOR2X1 XNOR2X1_80 ( .A(_abc_3927_n1649), .B(currentcol_15_), .Y(_abc_3927_n1650) );
	NOR2X1 NOR2X1_330 ( .A(_abc_3927_n1511), .B(_abc_3927_n1650), .Y(currentcol_15__FF_INPUT) );
	NAND2X1 NAND2X1_528 ( .A(currentrow_14_), .B(_abc_3927_n1586), .Y(_abc_3927_n1652) );
	XNOR2X1 XNOR2X1_81 ( .A(_abc_3927_n1652), .B(_abc_3927_n419), .Y(_abc_3927_n1653) );
	NOR2X1 NOR2X1_331 ( .A(_abc_3927_n1572), .B(_abc_3927_n1653), .Y(currentrow_15__FF_INPUT) );
	INVX1 INVX1_100 ( .A(reg_cr_value_15_), .Y(_abc_3927_n1655) );
	XNOR2X1 XNOR2X1_82 ( .A(currentrow_1_), .B(reg_ir_value_1_), .Y(_abc_3927_n1656) );
	XNOR2X1 XNOR2X1_83 ( .A(currentrow_0_), .B(reg_ir_value_0_), .Y(_abc_3927_n1657) );
	NAND2X1 NAND2X1_529 ( .A(_abc_3927_n1656), .B(_abc_3927_n1657), .Y(_abc_3927_n1658) );
	XNOR2X1 XNOR2X1_84 ( .A(currentrow_3_), .B(reg_ir_value_3_), .Y(_abc_3927_n1659) );
	XNOR2X1 XNOR2X1_85 ( .A(currentrow_2_), .B(reg_ir_value_2_), .Y(_abc_3927_n1660) );
	NAND2X1 NAND2X1_530 ( .A(_abc_3927_n1659), .B(_abc_3927_n1660), .Y(_abc_3927_n1661) );
	NOR2X1 NOR2X1_332 ( .A(_abc_3927_n1658), .B(_abc_3927_n1661), .Y(_abc_3927_n1662) );
	XNOR2X1 XNOR2X1_86 ( .A(currentrow_5_), .B(reg_ir_value_5_), .Y(_abc_3927_n1663) );
	XNOR2X1 XNOR2X1_87 ( .A(currentrow_4_), .B(reg_ir_value_4_), .Y(_abc_3927_n1664) );
	NAND2X1 NAND2X1_531 ( .A(_abc_3927_n1663), .B(_abc_3927_n1664), .Y(_abc_3927_n1665) );
	XNOR2X1 XNOR2X1_88 ( .A(currentrow_7_), .B(reg_ir_value_7_), .Y(_abc_3927_n1666) );
	XNOR2X1 XNOR2X1_89 ( .A(currentrow_6_), .B(reg_ir_value_6_), .Y(_abc_3927_n1667) );
	NAND2X1 NAND2X1_532 ( .A(_abc_3927_n1666), .B(_abc_3927_n1667), .Y(_abc_3927_n1668) );
	NOR2X1 NOR2X1_333 ( .A(_abc_3927_n1665), .B(_abc_3927_n1668), .Y(_abc_3927_n1669) );
	NAND2X1 NAND2X1_533 ( .A(_abc_3927_n1662), .B(_abc_3927_n1669), .Y(_abc_3927_n1670) );
	XNOR2X1 XNOR2X1_90 ( .A(currentrow_9_), .B(reg_ir_value_9_), .Y(_abc_3927_n1671) );
	XNOR2X1 XNOR2X1_91 ( .A(currentrow_8_), .B(reg_ir_value_8_), .Y(_abc_3927_n1672) );
	NAND2X1 NAND2X1_534 ( .A(_abc_3927_n1671), .B(_abc_3927_n1672), .Y(_abc_3927_n1673) );
	XNOR2X1 XNOR2X1_92 ( .A(currentrow_11_), .B(reg_ir_value_11_), .Y(_abc_3927_n1674) );
	XNOR2X1 XNOR2X1_93 ( .A(currentrow_10_), .B(reg_ir_value_10_), .Y(_abc_3927_n1675) );
	NAND2X1 NAND2X1_535 ( .A(_abc_3927_n1674), .B(_abc_3927_n1675), .Y(_abc_3927_n1676) );
	NOR2X1 NOR2X1_334 ( .A(_abc_3927_n1673), .B(_abc_3927_n1676), .Y(_abc_3927_n1677) );
	XNOR2X1 XNOR2X1_94 ( .A(currentrow_12_), .B(reg_ir_value_12_), .Y(_abc_3927_n1678) );
	XNOR2X1 XNOR2X1_95 ( .A(currentrow_13_), .B(reg_ir_value_13_), .Y(_abc_3927_n1679) );
	NAND2X1 NAND2X1_536 ( .A(_abc_3927_n1679), .B(_abc_3927_n1678), .Y(_abc_3927_n1680) );
	XNOR2X1 XNOR2X1_96 ( .A(currentrow_15_), .B(reg_ir_value_15_), .Y(_abc_3927_n1681) );
	XNOR2X1 XNOR2X1_97 ( .A(currentrow_14_), .B(reg_ir_value_14_), .Y(_abc_3927_n1682) );
	NAND2X1 NAND2X1_537 ( .A(_abc_3927_n1681), .B(_abc_3927_n1682), .Y(_abc_3927_n1683) );
	NOR2X1 NOR2X1_335 ( .A(_abc_3927_n1680), .B(_abc_3927_n1683), .Y(_abc_3927_n1684) );
	NAND2X1 NAND2X1_538 ( .A(_abc_3927_n1677), .B(_abc_3927_n1684), .Y(_abc_3927_n1685) );
	NOR2X1 NOR2X1_336 ( .A(_abc_3927_n1670), .B(_abc_3927_n1685), .Y(_abc_3927_n1686) );
	XNOR2X1 XNOR2X1_98 ( .A(currentcol_1_), .B(reg_ic_value_1_), .Y(_abc_3927_n1687) );
	XNOR2X1 XNOR2X1_99 ( .A(currentcol_0_), .B(reg_ic_value_0_), .Y(_abc_3927_n1688) );
	NAND2X1 NAND2X1_539 ( .A(_abc_3927_n1687), .B(_abc_3927_n1688), .Y(_abc_3927_n1689) );
	XNOR2X1 XNOR2X1_100 ( .A(currentcol_3_), .B(reg_ic_value_3_), .Y(_abc_3927_n1690) );
	XNOR2X1 XNOR2X1_101 ( .A(currentcol_2_), .B(reg_ic_value_2_), .Y(_abc_3927_n1691) );
	NAND2X1 NAND2X1_540 ( .A(_abc_3927_n1690), .B(_abc_3927_n1691), .Y(_abc_3927_n1692) );
	NOR2X1 NOR2X1_337 ( .A(_abc_3927_n1689), .B(_abc_3927_n1692), .Y(_abc_3927_n1693) );
	XNOR2X1 XNOR2X1_102 ( .A(currentcol_5_), .B(reg_ic_value_5_), .Y(_abc_3927_n1694) );
	XNOR2X1 XNOR2X1_103 ( .A(currentcol_4_), .B(reg_ic_value_4_), .Y(_abc_3927_n1695) );
	NAND2X1 NAND2X1_541 ( .A(_abc_3927_n1694), .B(_abc_3927_n1695), .Y(_abc_3927_n1696) );
	XNOR2X1 XNOR2X1_104 ( .A(currentcol_7_), .B(reg_ic_value_7_), .Y(_abc_3927_n1697) );
	XNOR2X1 XNOR2X1_105 ( .A(currentcol_6_), .B(reg_ic_value_6_), .Y(_abc_3927_n1698) );
	NAND2X1 NAND2X1_542 ( .A(_abc_3927_n1697), .B(_abc_3927_n1698), .Y(_abc_3927_n1699) );
	NOR2X1 NOR2X1_338 ( .A(_abc_3927_n1696), .B(_abc_3927_n1699), .Y(_abc_3927_n1700) );
	NAND2X1 NAND2X1_543 ( .A(_abc_3927_n1693), .B(_abc_3927_n1700), .Y(_abc_3927_n1701) );
	XNOR2X1 XNOR2X1_106 ( .A(currentcol_9_), .B(reg_ic_value_9_), .Y(_abc_3927_n1702) );
	XNOR2X1 XNOR2X1_107 ( .A(currentcol_8_), .B(reg_ic_value_8_), .Y(_abc_3927_n1703) );
	NAND2X1 NAND2X1_544 ( .A(_abc_3927_n1702), .B(_abc_3927_n1703), .Y(_abc_3927_n1704) );
	XNOR2X1 XNOR2X1_108 ( .A(currentcol_11_), .B(reg_ic_value_11_), .Y(_abc_3927_n1705) );
	XNOR2X1 XNOR2X1_109 ( .A(currentcol_10_), .B(reg_ic_value_10_), .Y(_abc_3927_n1706) );
	NAND2X1 NAND2X1_545 ( .A(_abc_3927_n1705), .B(_abc_3927_n1706), .Y(_abc_3927_n1707) );
	NOR2X1 NOR2X1_339 ( .A(_abc_3927_n1704), .B(_abc_3927_n1707), .Y(_abc_3927_n1708) );
	XNOR2X1 XNOR2X1_110 ( .A(currentcol_12_), .B(reg_ic_value_12_), .Y(_abc_3927_n1709) );
	XNOR2X1 XNOR2X1_111 ( .A(currentcol_13_), .B(reg_ic_value_13_), .Y(_abc_3927_n1710) );
	NAND2X1 NAND2X1_546 ( .A(_abc_3927_n1709), .B(_abc_3927_n1710), .Y(_abc_3927_n1711) );
	XNOR2X1 XNOR2X1_112 ( .A(currentcol_15_), .B(reg_ic_value_15_), .Y(_abc_3927_n1712) );
	XNOR2X1 XNOR2X1_113 ( .A(currentcol_14_), .B(reg_ic_value_14_), .Y(_abc_3927_n1713) );
	NAND2X1 NAND2X1_547 ( .A(_abc_3927_n1712), .B(_abc_3927_n1713), .Y(_abc_3927_n1714) );
	NOR2X1 NOR2X1_340 ( .A(_abc_3927_n1711), .B(_abc_3927_n1714), .Y(_abc_3927_n1715) );
	NAND2X1 NAND2X1_548 ( .A(_abc_3927_n1708), .B(_abc_3927_n1715), .Y(_abc_3927_n1716) );
	NOR2X1 NOR2X1_341 ( .A(_abc_3927_n1701), .B(_abc_3927_n1716), .Y(_abc_3927_n1717) );
	NAND2X1 NAND2X1_549 ( .A(_abc_3927_n1686), .B(_abc_3927_n1717), .Y(_abc_3927_n1718) );
	NOR2X1 NOR2X1_342 ( .A(_abc_3927_n1655), .B(_abc_3927_n1718), .Y(_abc_3927_n1719) );
	NOR2X1 NOR2X1_343 ( .A(_auto_iopadmap_cc_171_execute_5522), .B(_abc_3927_n1719), .Y(_abc_3927_n1720) );
	NAND2X1 NAND2X1_550 ( .A(addr_ir), .B(we), .Y(_abc_3927_n1721) );
	NAND2X1 NAND2X1_551 ( .A(_abc_3927_n365), .B(_abc_3927_n1721), .Y(_abc_3927_n1722) );
	NOR2X1 NOR2X1_344 ( .A(_abc_3927_n1722), .B(_abc_3927_n1720), .Y(irq_FF_INPUT) );
	NOR2X1 NOR2X1_345 ( .A(reg_cr_value_0_), .B(_abc_3927_n815_1), .Y(_auto_iopadmap_cc_171_execute_5516) );
	AND2X2 AND2X2_117 ( .A(_abc_3927_n419), .B(reg_vb_value_15_), .Y(_abc_3927_n1725) );
	NOR2X1 NOR2X1_346 ( .A(reg_vb_value_15_), .B(_abc_3927_n419), .Y(_abc_3927_n1726) );
	NOR2X1 NOR2X1_347 ( .A(_abc_3927_n1726), .B(_abc_3927_n1725), .Y(_abc_3927_n1727) );
	AND2X2 AND2X2_118 ( .A(_abc_3927_n423), .B(reg_vb_value_14_), .Y(_abc_3927_n1728) );
	NOR2X1 NOR2X1_348 ( .A(reg_vb_value_14_), .B(_abc_3927_n423), .Y(_abc_3927_n1729) );
	NOR2X1 NOR2X1_349 ( .A(_abc_3927_n1729), .B(_abc_3927_n1728), .Y(_abc_3927_n1730) );
	NAND2X1 NAND2X1_552 ( .A(_abc_3927_n1727), .B(_abc_3927_n1730), .Y(_abc_3927_n1731) );
	INVX1 INVX1_101 ( .A(_abc_3927_n1731), .Y(_abc_3927_n1732) );
	XOR2X1 XOR2X1_38 ( .A(reg_vb_value_13_), .B(currentrow_13_), .Y(_abc_3927_n1733) );
	XOR2X1 XOR2X1_39 ( .A(reg_vb_value_12_), .B(currentrow_12_), .Y(_abc_3927_n1734) );
	NOR2X1 NOR2X1_350 ( .A(_abc_3927_n1733), .B(_abc_3927_n1734), .Y(_abc_3927_n1735) );
	NAND2X1 NAND2X1_553 ( .A(_abc_3927_n1735), .B(_abc_3927_n1732), .Y(_abc_3927_n1736) );
	NAND2X1 NAND2X1_554 ( .A(reg_vb_value_11_), .B(_abc_3927_n438_1), .Y(_abc_3927_n1737) );
	OR2X2 OR2X2_66 ( .A(_abc_3927_n438_1), .B(reg_vb_value_11_), .Y(_abc_3927_n1738) );
	NAND2X1 NAND2X1_555 ( .A(_abc_3927_n1737), .B(_abc_3927_n1738), .Y(_abc_3927_n1739) );
	XOR2X1 XOR2X1_40 ( .A(reg_vb_value_10_), .B(currentrow_10_), .Y(_abc_3927_n1740) );
	NOR2X1 NOR2X1_351 ( .A(_abc_3927_n1740), .B(_abc_3927_n1739), .Y(_abc_3927_n1741) );
	INVX1 INVX1_102 ( .A(reg_vb_value_8_), .Y(_abc_3927_n1742) );
	NAND2X1 NAND2X1_556 ( .A(currentrow_8_), .B(_abc_3927_n1742), .Y(_abc_3927_n1743) );
	OR2X2 OR2X2_67 ( .A(_abc_3927_n446), .B(reg_vb_value_9_), .Y(_abc_3927_n1744) );
	NAND2X1 NAND2X1_557 ( .A(_abc_3927_n1743), .B(_abc_3927_n1744), .Y(_abc_3927_n1745) );
	NAND2X1 NAND2X1_558 ( .A(reg_vb_value_9_), .B(_abc_3927_n446), .Y(_abc_3927_n1746) );
	NOR2X1 NOR2X1_352 ( .A(currentrow_8_), .B(_abc_3927_n1742), .Y(_abc_3927_n1747) );
	INVX1 INVX1_103 ( .A(_abc_3927_n1747), .Y(_abc_3927_n1748) );
	NAND2X1 NAND2X1_559 ( .A(_abc_3927_n1746), .B(_abc_3927_n1748), .Y(_abc_3927_n1749) );
	NOR2X1 NOR2X1_353 ( .A(_abc_3927_n1745), .B(_abc_3927_n1749), .Y(_abc_3927_n1750) );
	NAND2X1 NAND2X1_560 ( .A(_abc_3927_n1741), .B(_abc_3927_n1750), .Y(_abc_3927_n1751) );
	NOR2X1 NOR2X1_354 ( .A(_abc_3927_n1751), .B(_abc_3927_n1736), .Y(_abc_3927_n1752) );
	NOR2X1 NOR2X1_355 ( .A(reg_vb_value_7_), .B(_abc_3927_n456), .Y(_abc_3927_n1753) );
	NAND2X1 NAND2X1_561 ( .A(reg_vb_value_7_), .B(_abc_3927_n456), .Y(_abc_3927_n1754) );
	INVX1 INVX1_104 ( .A(_abc_3927_n1754), .Y(_abc_3927_n1755) );
	NOR2X1 NOR2X1_356 ( .A(_abc_3927_n1753), .B(_abc_3927_n1755), .Y(_abc_3927_n1756) );
	XNOR2X1 XNOR2X1_114 ( .A(reg_vb_value_6_), .B(currentrow_6_), .Y(_abc_3927_n1757) );
	AND2X2 AND2X2_119 ( .A(_abc_3927_n1756), .B(_abc_3927_n1757), .Y(_abc_3927_n1758) );
	OR2X2 OR2X2_68 ( .A(_abc_3927_n462), .B(reg_vb_value_5_), .Y(_abc_3927_n1759) );
	INVX1 INVX1_105 ( .A(reg_vb_value_4_), .Y(_abc_3927_n1760) );
	NAND2X1 NAND2X1_562 ( .A(currentrow_4_), .B(_abc_3927_n1760), .Y(_abc_3927_n1761) );
	NAND2X1 NAND2X1_563 ( .A(_abc_3927_n1761), .B(_abc_3927_n1759), .Y(_abc_3927_n1762) );
	NOR2X1 NOR2X1_357 ( .A(currentrow_4_), .B(_abc_3927_n1760), .Y(_abc_3927_n1763) );
	INVX1 INVX1_106 ( .A(_abc_3927_n1763), .Y(_abc_3927_n1764) );
	NAND2X1 NAND2X1_564 ( .A(reg_vb_value_5_), .B(_abc_3927_n462), .Y(_abc_3927_n1765) );
	NAND2X1 NAND2X1_565 ( .A(_abc_3927_n1765), .B(_abc_3927_n1764), .Y(_abc_3927_n1766) );
	NOR2X1 NOR2X1_358 ( .A(_abc_3927_n1762), .B(_abc_3927_n1766), .Y(_abc_3927_n1767) );
	NAND2X1 NAND2X1_566 ( .A(_abc_3927_n1767), .B(_abc_3927_n1758), .Y(_abc_3927_n1768) );
	NAND2X1 NAND2X1_567 ( .A(reg_vb_value_3_), .B(_abc_3927_n472), .Y(_abc_3927_n1769) );
	OR2X2 OR2X2_69 ( .A(_abc_3927_n472), .B(reg_vb_value_3_), .Y(_abc_3927_n1770) );
	NAND2X1 NAND2X1_568 ( .A(_abc_3927_n1769), .B(_abc_3927_n1770), .Y(_abc_3927_n1771) );
	XOR2X1 XOR2X1_41 ( .A(reg_vb_value_2_), .B(currentrow_2_), .Y(_abc_3927_n1772) );
	NOR2X1 NOR2X1_359 ( .A(_abc_3927_n1772), .B(_abc_3927_n1771), .Y(_abc_3927_n1773) );
	INVX1 INVX1_107 ( .A(reg_vb_value_0_), .Y(_abc_3927_n1774) );
	NOR2X1 NOR2X1_360 ( .A(currentrow_0_), .B(_abc_3927_n1774), .Y(_abc_3927_n1775) );
	NAND2X1 NAND2X1_569 ( .A(currentrow_0_), .B(_abc_3927_n1774), .Y(_abc_3927_n1776) );
	XNOR2X1 XNOR2X1_115 ( .A(reg_vb_value_1_), .B(currentrow_1_), .Y(_abc_3927_n1777) );
	NAND2X1 NAND2X1_570 ( .A(_abc_3927_n1776), .B(_abc_3927_n1777), .Y(_abc_3927_n1778) );
	NOR2X1 NOR2X1_361 ( .A(_abc_3927_n1775), .B(_abc_3927_n1778), .Y(_abc_3927_n1779) );
	NAND2X1 NAND2X1_571 ( .A(_abc_3927_n1773), .B(_abc_3927_n1779), .Y(_abc_3927_n1780) );
	NOR2X1 NOR2X1_362 ( .A(_abc_3927_n1780), .B(_abc_3927_n1768), .Y(_abc_3927_n1781) );
	NAND2X1 NAND2X1_572 ( .A(_abc_3927_n1781), .B(_abc_3927_n1752), .Y(_abc_3927_n1782) );
	INVX1 INVX1_108 ( .A(_abc_3927_n1768), .Y(_abc_3927_n1783) );
	NAND2X1 NAND2X1_573 ( .A(reg_vb_value_1_), .B(_abc_3927_n478_1), .Y(_abc_3927_n1784) );
	NAND2X1 NAND2X1_574 ( .A(_abc_3927_n1784), .B(_abc_3927_n1778), .Y(_abc_3927_n1785) );
	NAND2X1 NAND2X1_575 ( .A(_abc_3927_n1773), .B(_abc_3927_n1785), .Y(_abc_3927_n1786) );
	AND2X2 AND2X2_120 ( .A(_abc_3927_n486_1), .B(reg_vb_value_2_), .Y(_abc_3927_n1787) );
	NAND2X1 NAND2X1_576 ( .A(_abc_3927_n1787), .B(_abc_3927_n1770), .Y(_abc_3927_n1788) );
	AND2X2 AND2X2_121 ( .A(_abc_3927_n1788), .B(_abc_3927_n1769), .Y(_abc_3927_n1789) );
	NAND2X1 NAND2X1_577 ( .A(_abc_3927_n1789), .B(_abc_3927_n1786), .Y(_abc_3927_n1790) );
	NAND2X1 NAND2X1_578 ( .A(_abc_3927_n1790), .B(_abc_3927_n1783), .Y(_abc_3927_n1791) );
	NAND2X1 NAND2X1_579 ( .A(_abc_3927_n1763), .B(_abc_3927_n1759), .Y(_abc_3927_n1792) );
	NAND2X1 NAND2X1_580 ( .A(_abc_3927_n1765), .B(_abc_3927_n1792), .Y(_abc_3927_n1793) );
	NAND2X1 NAND2X1_581 ( .A(_abc_3927_n1793), .B(_abc_3927_n1758), .Y(_abc_3927_n1794) );
	NAND2X1 NAND2X1_582 ( .A(reg_vb_value_6_), .B(_abc_3927_n496), .Y(_abc_3927_n1795) );
	NOR2X1 NOR2X1_363 ( .A(_abc_3927_n1795), .B(_abc_3927_n1753), .Y(_abc_3927_n1796) );
	NOR2X1 NOR2X1_364 ( .A(_abc_3927_n1755), .B(_abc_3927_n1796), .Y(_abc_3927_n1797) );
	AND2X2 AND2X2_122 ( .A(_abc_3927_n1794), .B(_abc_3927_n1797), .Y(_abc_3927_n1798) );
	NAND2X1 NAND2X1_583 ( .A(_abc_3927_n1798), .B(_abc_3927_n1791), .Y(_abc_3927_n1799) );
	NAND2X1 NAND2X1_584 ( .A(_abc_3927_n1752), .B(_abc_3927_n1799), .Y(_abc_3927_n1800) );
	NAND2X1 NAND2X1_585 ( .A(_abc_3927_n1747), .B(_abc_3927_n1744), .Y(_abc_3927_n1801) );
	NAND2X1 NAND2X1_586 ( .A(_abc_3927_n1746), .B(_abc_3927_n1801), .Y(_abc_3927_n1802) );
	NAND2X1 NAND2X1_587 ( .A(_abc_3927_n1802), .B(_abc_3927_n1741), .Y(_abc_3927_n1803) );
	AND2X2 AND2X2_123 ( .A(_abc_3927_n506), .B(reg_vb_value_10_), .Y(_abc_3927_n1804) );
	NAND2X1 NAND2X1_588 ( .A(_abc_3927_n1804), .B(_abc_3927_n1738), .Y(_abc_3927_n1805) );
	AND2X2 AND2X2_124 ( .A(_abc_3927_n1805), .B(_abc_3927_n1737), .Y(_abc_3927_n1806) );
	AND2X2 AND2X2_125 ( .A(_abc_3927_n1803), .B(_abc_3927_n1806), .Y(_abc_3927_n1807) );
	NOR2X1 NOR2X1_365 ( .A(_abc_3927_n1736), .B(_abc_3927_n1807), .Y(_abc_3927_n1808) );
	NAND2X1 NAND2X1_589 ( .A(reg_vb_value_13_), .B(_abc_3927_n432_1), .Y(_abc_3927_n1809) );
	NAND2X1 NAND2X1_590 ( .A(reg_vb_value_12_), .B(_abc_3927_n428_1), .Y(_abc_3927_n1810) );
	OR2X2 OR2X2_70 ( .A(_abc_3927_n1733), .B(_abc_3927_n1810), .Y(_abc_3927_n1811) );
	NAND2X1 NAND2X1_591 ( .A(_abc_3927_n1809), .B(_abc_3927_n1811), .Y(_abc_3927_n1812) );
	NAND2X1 NAND2X1_592 ( .A(_abc_3927_n1812), .B(_abc_3927_n1732), .Y(_abc_3927_n1813) );
	AND2X2 AND2X2_126 ( .A(_abc_3927_n1727), .B(_abc_3927_n1728), .Y(_abc_3927_n1814) );
	NOR2X1 NOR2X1_366 ( .A(_abc_3927_n1725), .B(_abc_3927_n1814), .Y(_abc_3927_n1815) );
	NAND2X1 NAND2X1_593 ( .A(_abc_3927_n1815), .B(_abc_3927_n1813), .Y(_abc_3927_n1816) );
	NOR2X1 NOR2X1_367 ( .A(_abc_3927_n1816), .B(_abc_3927_n1808), .Y(_abc_3927_n1817) );
	NAND2X1 NAND2X1_594 ( .A(_abc_3927_n1817), .B(_abc_3927_n1800), .Y(_abc_3927_n1818) );
	NAND2X1 NAND2X1_595 ( .A(_abc_3927_n1782), .B(_abc_3927_n1818), .Y(_abc_3927_n1819) );
	XNOR2X1 XNOR2X1_116 ( .A(_abc_3927_n1819), .B(reg_cr_value_13_), .Y(_abc_3927_n1528) );
	NOR2X1 NOR2X1_368 ( .A(reg_hb_value_14_), .B(_abc_3927_n524), .Y(_abc_3927_n1821) );
	NOR2X1 NOR2X1_369 ( .A(reg_hb_value_15_), .B(_abc_3927_n520), .Y(_abc_3927_n1822) );
	INVX1 INVX1_109 ( .A(_abc_3927_n1822), .Y(_abc_3927_n1823) );
	NAND2X1 NAND2X1_596 ( .A(reg_hb_value_15_), .B(_abc_3927_n520), .Y(_abc_3927_n1824) );
	NAND2X1 NAND2X1_597 ( .A(_abc_3927_n1824), .B(_abc_3927_n1823), .Y(_abc_3927_n1825) );
	NAND2X1 NAND2X1_598 ( .A(reg_hb_value_14_), .B(_abc_3927_n524), .Y(_abc_3927_n1826) );
	INVX1 INVX1_110 ( .A(_abc_3927_n1826), .Y(_abc_3927_n1827) );
	OR2X2 OR2X2_71 ( .A(_abc_3927_n1825), .B(_abc_3927_n1827), .Y(_abc_3927_n1828) );
	NOR2X1 NOR2X1_370 ( .A(_abc_3927_n1821), .B(_abc_3927_n1828), .Y(_abc_3927_n1829) );
	NAND2X1 NAND2X1_599 ( .A(reg_hb_value_13_), .B(_abc_3927_n529), .Y(_abc_3927_n1830) );
	NAND2X1 NAND2X1_600 ( .A(reg_hb_value_12_), .B(_abc_3927_n531), .Y(_abc_3927_n1831) );
	NAND2X1 NAND2X1_601 ( .A(_abc_3927_n1830), .B(_abc_3927_n1831), .Y(_abc_3927_n1832) );
	OR2X2 OR2X2_72 ( .A(_abc_3927_n529), .B(reg_hb_value_13_), .Y(_abc_3927_n1833) );
	OR2X2 OR2X2_73 ( .A(_abc_3927_n531), .B(reg_hb_value_12_), .Y(_abc_3927_n1834) );
	NAND2X1 NAND2X1_602 ( .A(_abc_3927_n1833), .B(_abc_3927_n1834), .Y(_abc_3927_n1835) );
	NOR2X1 NOR2X1_371 ( .A(_abc_3927_n1832), .B(_abc_3927_n1835), .Y(_abc_3927_n1836) );
	NAND2X1 NAND2X1_603 ( .A(_abc_3927_n1836), .B(_abc_3927_n1829), .Y(_abc_3927_n1837) );
	NAND2X1 NAND2X1_604 ( .A(reg_hb_value_11_), .B(_abc_3927_n539), .Y(_abc_3927_n1838) );
	NAND2X1 NAND2X1_605 ( .A(reg_hb_value_10_), .B(_abc_3927_n604), .Y(_abc_3927_n1839) );
	NAND2X1 NAND2X1_606 ( .A(_abc_3927_n1838), .B(_abc_3927_n1839), .Y(_abc_3927_n1840) );
	OR2X2 OR2X2_74 ( .A(_abc_3927_n539), .B(reg_hb_value_11_), .Y(_abc_3927_n1841) );
	OR2X2 OR2X2_75 ( .A(_abc_3927_n604), .B(reg_hb_value_10_), .Y(_abc_3927_n1842) );
	NAND2X1 NAND2X1_607 ( .A(_abc_3927_n1841), .B(_abc_3927_n1842), .Y(_abc_3927_n1843) );
	NOR2X1 NOR2X1_372 ( .A(_abc_3927_n1840), .B(_abc_3927_n1843), .Y(_abc_3927_n1844) );
	NAND2X1 NAND2X1_608 ( .A(reg_hb_value_9_), .B(_abc_3927_n546), .Y(_abc_3927_n1845) );
	NAND2X1 NAND2X1_609 ( .A(reg_hb_value_8_), .B(_abc_3927_n548), .Y(_abc_3927_n1846) );
	NAND2X1 NAND2X1_610 ( .A(_abc_3927_n1845), .B(_abc_3927_n1846), .Y(_abc_3927_n1847) );
	OR2X2 OR2X2_76 ( .A(_abc_3927_n546), .B(reg_hb_value_9_), .Y(_abc_3927_n1848) );
	OR2X2 OR2X2_77 ( .A(_abc_3927_n548), .B(reg_hb_value_8_), .Y(_abc_3927_n1849) );
	NAND2X1 NAND2X1_611 ( .A(_abc_3927_n1848), .B(_abc_3927_n1849), .Y(_abc_3927_n1850) );
	NOR2X1 NOR2X1_373 ( .A(_abc_3927_n1847), .B(_abc_3927_n1850), .Y(_abc_3927_n1851) );
	NAND2X1 NAND2X1_612 ( .A(_abc_3927_n1851), .B(_abc_3927_n1844), .Y(_abc_3927_n1852) );
	NOR2X1 NOR2X1_374 ( .A(_abc_3927_n1852), .B(_abc_3927_n1837), .Y(_abc_3927_n1853) );
	NOR2X1 NOR2X1_375 ( .A(reg_hb_value_6_), .B(_abc_3927_n562), .Y(_abc_3927_n1854) );
	NOR2X1 NOR2X1_376 ( .A(reg_hb_value_7_), .B(_abc_3927_n663), .Y(_abc_3927_n1855) );
	INVX1 INVX1_111 ( .A(_abc_3927_n1855), .Y(_abc_3927_n1856) );
	NAND2X1 NAND2X1_613 ( .A(reg_hb_value_7_), .B(_abc_3927_n663), .Y(_abc_3927_n1857) );
	NAND2X1 NAND2X1_614 ( .A(_abc_3927_n1857), .B(_abc_3927_n1856), .Y(_abc_3927_n1858) );
	NAND2X1 NAND2X1_615 ( .A(reg_hb_value_6_), .B(_abc_3927_n562), .Y(_abc_3927_n1859) );
	INVX1 INVX1_112 ( .A(_abc_3927_n1859), .Y(_abc_3927_n1860) );
	OR2X2 OR2X2_78 ( .A(_abc_3927_n1858), .B(_abc_3927_n1860), .Y(_abc_3927_n1861) );
	NOR2X1 NOR2X1_377 ( .A(_abc_3927_n1854), .B(_abc_3927_n1861), .Y(_abc_3927_n1862) );
	NAND2X1 NAND2X1_616 ( .A(reg_hb_value_5_), .B(_abc_3927_n567), .Y(_abc_3927_n1863) );
	NAND2X1 NAND2X1_617 ( .A(reg_hb_value_4_), .B(_abc_3927_n569), .Y(_abc_3927_n1864) );
	NAND2X1 NAND2X1_618 ( .A(_abc_3927_n1863), .B(_abc_3927_n1864), .Y(_abc_3927_n1865) );
	OR2X2 OR2X2_79 ( .A(_abc_3927_n567), .B(reg_hb_value_5_), .Y(_abc_3927_n1866) );
	OR2X2 OR2X2_80 ( .A(_abc_3927_n569), .B(reg_hb_value_4_), .Y(_abc_3927_n1867) );
	NAND2X1 NAND2X1_619 ( .A(_abc_3927_n1866), .B(_abc_3927_n1867), .Y(_abc_3927_n1868) );
	NOR2X1 NOR2X1_378 ( .A(_abc_3927_n1865), .B(_abc_3927_n1868), .Y(_abc_3927_n1869) );
	NAND2X1 NAND2X1_620 ( .A(_abc_3927_n1869), .B(_abc_3927_n1862), .Y(_abc_3927_n1870) );
	NAND2X1 NAND2X1_621 ( .A(reg_hb_value_3_), .B(_abc_3927_n577), .Y(_abc_3927_n1871) );
	OR2X2 OR2X2_81 ( .A(_abc_3927_n577), .B(reg_hb_value_3_), .Y(_abc_3927_n1872) );
	NAND2X1 NAND2X1_622 ( .A(_abc_3927_n1871), .B(_abc_3927_n1872), .Y(_abc_3927_n1873) );
	XOR2X1 XOR2X1_42 ( .A(currentcol_2_), .B(reg_hb_value_2_), .Y(_abc_3927_n1874) );
	NOR2X1 NOR2X1_379 ( .A(_abc_3927_n1874), .B(_abc_3927_n1873), .Y(_abc_3927_n1875) );
	INVX1 INVX1_113 ( .A(reg_hb_value_1_), .Y(_abc_3927_n1876) );
	NOR2X1 NOR2X1_380 ( .A(currentcol_1_), .B(_abc_3927_n1876), .Y(_abc_3927_n1877) );
	INVX1 INVX1_114 ( .A(_abc_3927_n1877), .Y(_abc_3927_n1878) );
	OR2X2 OR2X2_82 ( .A(_abc_3927_n585), .B(reg_hb_value_0_), .Y(_abc_3927_n1879) );
	NOR2X1 NOR2X1_381 ( .A(reg_hb_value_1_), .B(_abc_3927_n583), .Y(_abc_3927_n1880) );
	NOR2X1 NOR2X1_382 ( .A(_abc_3927_n1877), .B(_abc_3927_n1880), .Y(_abc_3927_n1881) );
	NAND2X1 NAND2X1_623 ( .A(_abc_3927_n1879), .B(_abc_3927_n1881), .Y(_abc_3927_n1882) );
	NAND2X1 NAND2X1_624 ( .A(_abc_3927_n1878), .B(_abc_3927_n1882), .Y(_abc_3927_n1883) );
	NAND2X1 NAND2X1_625 ( .A(_abc_3927_n1875), .B(_abc_3927_n1883), .Y(_abc_3927_n1884) );
	AND2X2 AND2X2_127 ( .A(_abc_3927_n591), .B(reg_hb_value_2_), .Y(_abc_3927_n1885) );
	NAND2X1 NAND2X1_626 ( .A(_abc_3927_n1885), .B(_abc_3927_n1872), .Y(_abc_3927_n1886) );
	AND2X2 AND2X2_128 ( .A(_abc_3927_n1886), .B(_abc_3927_n1871), .Y(_abc_3927_n1887) );
	AND2X2 AND2X2_129 ( .A(_abc_3927_n1884), .B(_abc_3927_n1887), .Y(_abc_3927_n1888) );
	OR2X2 OR2X2_83 ( .A(_abc_3927_n1888), .B(_abc_3927_n1870), .Y(_abc_3927_n1889) );
	NAND2X1 NAND2X1_627 ( .A(_abc_3927_n1860), .B(_abc_3927_n1856), .Y(_abc_3927_n1890) );
	NAND2X1 NAND2X1_628 ( .A(_abc_3927_n1857), .B(_abc_3927_n1890), .Y(_abc_3927_n1891) );
	AND2X2 AND2X2_130 ( .A(_abc_3927_n1865), .B(_abc_3927_n1866), .Y(_abc_3927_n1892) );
	AND2X2 AND2X2_131 ( .A(_abc_3927_n1862), .B(_abc_3927_n1892), .Y(_abc_3927_n1893) );
	NOR2X1 NOR2X1_383 ( .A(_abc_3927_n1891), .B(_abc_3927_n1893), .Y(_abc_3927_n1894) );
	NAND2X1 NAND2X1_629 ( .A(_abc_3927_n1894), .B(_abc_3927_n1889), .Y(_abc_3927_n1895) );
	NAND2X1 NAND2X1_630 ( .A(_abc_3927_n1853), .B(_abc_3927_n1895), .Y(_abc_3927_n1896) );
	NAND2X1 NAND2X1_631 ( .A(_abc_3927_n1841), .B(_abc_3927_n1840), .Y(_abc_3927_n1897) );
	AND2X2 AND2X2_132 ( .A(_abc_3927_n1847), .B(_abc_3927_n1848), .Y(_abc_3927_n1898) );
	NAND2X1 NAND2X1_632 ( .A(_abc_3927_n1898), .B(_abc_3927_n1844), .Y(_abc_3927_n1899) );
	AND2X2 AND2X2_133 ( .A(_abc_3927_n1899), .B(_abc_3927_n1897), .Y(_abc_3927_n1900) );
	NOR2X1 NOR2X1_384 ( .A(_abc_3927_n1900), .B(_abc_3927_n1837), .Y(_abc_3927_n1901) );
	AND2X2 AND2X2_134 ( .A(_abc_3927_n1832), .B(_abc_3927_n1833), .Y(_abc_3927_n1902) );
	NAND2X1 NAND2X1_633 ( .A(_abc_3927_n1902), .B(_abc_3927_n1829), .Y(_abc_3927_n1903) );
	NAND2X1 NAND2X1_634 ( .A(_abc_3927_n1827), .B(_abc_3927_n1823), .Y(_abc_3927_n1904) );
	AND2X2 AND2X2_135 ( .A(_abc_3927_n1904), .B(_abc_3927_n1824), .Y(_abc_3927_n1905) );
	NAND2X1 NAND2X1_635 ( .A(_abc_3927_n1905), .B(_abc_3927_n1903), .Y(_abc_3927_n1906) );
	NOR2X1 NOR2X1_385 ( .A(_abc_3927_n1906), .B(_abc_3927_n1901), .Y(_abc_3927_n1907) );
	NAND2X1 NAND2X1_636 ( .A(_abc_3927_n1907), .B(_abc_3927_n1896), .Y(_abc_3927_n1908) );
	NAND2X1 NAND2X1_637 ( .A(reg_hb_value_0_), .B(_abc_3927_n585), .Y(_abc_3927_n1909) );
	NAND2X1 NAND2X1_638 ( .A(_abc_3927_n1909), .B(_abc_3927_n1875), .Y(_abc_3927_n1910) );
	OR2X2 OR2X2_84 ( .A(_abc_3927_n1910), .B(_abc_3927_n1882), .Y(_abc_3927_n1911) );
	NOR2X1 NOR2X1_386 ( .A(_abc_3927_n1911), .B(_abc_3927_n1870), .Y(_abc_3927_n1912) );
	NAND2X1 NAND2X1_639 ( .A(_abc_3927_n1853), .B(_abc_3927_n1912), .Y(_abc_3927_n1913) );
	NAND2X1 NAND2X1_640 ( .A(_abc_3927_n1913), .B(_abc_3927_n1908), .Y(_abc_3927_n1914) );
	XNOR2X1 XNOR2X1_117 ( .A(_abc_3927_n1914), .B(reg_cr_value_14_), .Y(_abc_3927_n1531) );
	BUFX2 BUFX2_1 ( .A(currentaddr_0_), .Y(pixaddr[0]) );
	BUFX2 BUFX2_2 ( .A(currentaddr_1_), .Y(pixaddr[1]) );
	BUFX2 BUFX2_3 ( .A(currentaddr_2_), .Y(pixaddr[2]) );
	BUFX2 BUFX2_4 ( .A(currentaddr_3_), .Y(pixaddr[3]) );
	BUFX2 BUFX2_5 ( .A(currentaddr_4_), .Y(pixaddr[4]) );
	BUFX2 BUFX2_6 ( .A(currentaddr_5_), .Y(pixaddr[5]) );
	BUFX2 BUFX2_7 ( .A(currentaddr_6_), .Y(pixaddr[6]) );
	BUFX2 BUFX2_8 ( .A(currentaddr_7_), .Y(pixaddr[7]) );
	BUFX2 BUFX2_9 ( .A(currentaddr_8_), .Y(pixaddr[8]) );
	BUFX2 BUFX2_10 ( .A(currentaddr_9_), .Y(pixaddr[9]) );
	BUFX2 BUFX2_11 ( .A(currentaddr_10_), .Y(pixaddr[10]) );
	BUFX2 BUFX2_12 ( .A(currentaddr_11_), .Y(pixaddr[11]) );
	BUFX2 BUFX2_13 ( .A(currentaddr_12_), .Y(pixaddr[12]) );
	BUFX2 BUFX2_14 ( .A(currentaddr_13_), .Y(pixaddr[13]) );
	BUFX2 BUFX2_15 ( .A(currentaddr_14_), .Y(pixaddr[14]) );
	BUFX2 BUFX2_16 ( .A(currentaddr_15_), .Y(pixaddr[15]) );
	BUFX2 BUFX2_17 ( .A(currentaddr_16_), .Y(pixaddr[16]) );
	BUFX2 BUFX2_18 ( .A(currentaddr_17_), .Y(pixaddr[17]) );
	BUFX2 BUFX2_19 ( .A(currentaddr_18_), .Y(pixaddr[18]) );
	BUFX2 BUFX2_20 ( .A(currentaddr_19_), .Y(pixaddr[19]) );
	BUFX2 BUFX2_21 ( .A(currentaddr_20_), .Y(pixaddr[20]) );
	BUFX2 BUFX2_22 ( .A(currentaddr_21_), .Y(pixaddr[21]) );
	BUFX2 BUFX2_23 ( .A(currentaddr_22_), .Y(pixaddr[22]) );
	BUFX2 BUFX2_24 ( .A(currentaddr_23_), .Y(pixaddr[23]) );
	BUFX2 BUFX2_25 ( .A(currentaddr_24_), .Y(pixaddr[24]) );
	BUFX2 BUFX2_26 ( .A(currentaddr_25_), .Y(pixaddr[25]) );
	BUFX2 BUFX2_27 ( .A(currentaddr_26_), .Y(pixaddr[26]) );
	BUFX2 BUFX2_28 ( .A(currentaddr_27_), .Y(pixaddr[27]) );
	BUFX2 BUFX2_29 ( .A(currentaddr_28_), .Y(pixaddr[28]) );
	BUFX2 BUFX2_30 ( .A(currentaddr_29_), .Y(pixaddr[29]) );
	BUFX2 BUFX2_31 ( .A(currentaddr_30_), .Y(pixaddr[30]) );
	BUFX2 BUFX2_32 ( .A(currentaddr_31_), .Y(pixaddr[31]) );
	BUFX2 BUFX2_33 ( .A(reg_cr_value_5_), .Y(clksel[0]) );
	BUFX2 BUFX2_34 ( .A(reg_cr_value_6_), .Y(clksel[1]) );
	BUFX2 BUFX2_35 ( .A(reg_cr_value_7_), .Y(clksel[2]) );
	BUFX2 BUFX2_36 ( .A(_auto_iopadmap_cc_171_execute_5516), .Y(ven) );
	BUFX2 BUFX2_37 ( .A(_abc_3927_n1531), .Y(hs) );
	BUFX2 BUFX2_38 ( .A(_abc_3927_n1528), .Y(vs) );
	BUFX2 BUFX2_39 ( .A(_auto_iopadmap_cc_171_execute_5522), .Y(irq) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(irq_FF_INPUT), .Q(_auto_iopadmap_cc_171_execute_5522) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(currentrow_0__FF_INPUT), .Q(currentrow_0_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(currentrow_1__FF_INPUT), .Q(currentrow_1_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(currentrow_2__FF_INPUT), .Q(currentrow_2_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(currentrow_3__FF_INPUT), .Q(currentrow_3_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(currentrow_4__FF_INPUT), .Q(currentrow_4_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(currentrow_5__FF_INPUT), .Q(currentrow_5_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(currentrow_6__FF_INPUT), .Q(currentrow_6_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(currentrow_7__FF_INPUT), .Q(currentrow_7_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(currentrow_8__FF_INPUT), .Q(currentrow_8_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(currentrow_9__FF_INPUT), .Q(currentrow_9_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(currentrow_10__FF_INPUT), .Q(currentrow_10_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(currentrow_11__FF_INPUT), .Q(currentrow_11_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(currentrow_12__FF_INPUT), .Q(currentrow_12_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(currentrow_13__FF_INPUT), .Q(currentrow_13_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(currentrow_14__FF_INPUT), .Q(currentrow_14_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(currentrow_15__FF_INPUT), .Q(currentrow_15_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(currentcol_0__FF_INPUT), .Q(currentcol_0_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(currentcol_1__FF_INPUT), .Q(currentcol_1_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(currentcol_2__FF_INPUT), .Q(currentcol_2_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(currentcol_3__FF_INPUT), .Q(currentcol_3_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(currentcol_4__FF_INPUT), .Q(currentcol_4_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(currentcol_5__FF_INPUT), .Q(currentcol_5_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(currentcol_6__FF_INPUT), .Q(currentcol_6_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(currentcol_7__FF_INPUT), .Q(currentcol_7_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(currentcol_8__FF_INPUT), .Q(currentcol_8_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(currentcol_9__FF_INPUT), .Q(currentcol_9_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(currentcol_10__FF_INPUT), .Q(currentcol_10_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(currentcol_11__FF_INPUT), .Q(currentcol_11_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(currentcol_12__FF_INPUT), .Q(currentcol_12_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(currentcol_13__FF_INPUT), .Q(currentcol_13_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(currentcol_14__FF_INPUT), .Q(currentcol_14_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(currentcol_15__FF_INPUT), .Q(currentcol_15_) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(currentaddr_0__FF_INPUT), .Q(currentaddr_0_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(currentaddr_1__FF_INPUT), .Q(currentaddr_1_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(currentaddr_2__FF_INPUT), .Q(currentaddr_2_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(currentaddr_3__FF_INPUT), .Q(currentaddr_3_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(currentaddr_4__FF_INPUT), .Q(currentaddr_4_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(currentaddr_5__FF_INPUT), .Q(currentaddr_5_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(currentaddr_6__FF_INPUT), .Q(currentaddr_6_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(currentaddr_7__FF_INPUT), .Q(currentaddr_7_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(currentaddr_8__FF_INPUT), .Q(currentaddr_8_) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(currentaddr_9__FF_INPUT), .Q(currentaddr_9_) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(currentaddr_10__FF_INPUT), .Q(currentaddr_10_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(currentaddr_11__FF_INPUT), .Q(currentaddr_11_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(currentaddr_12__FF_INPUT), .Q(currentaddr_12_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(currentaddr_13__FF_INPUT), .Q(currentaddr_13_) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(currentaddr_14__FF_INPUT), .Q(currentaddr_14_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(currentaddr_15__FF_INPUT), .Q(currentaddr_15_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(currentaddr_16__FF_INPUT), .Q(currentaddr_16_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(currentaddr_17__FF_INPUT), .Q(currentaddr_17_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(currentaddr_18__FF_INPUT), .Q(currentaddr_18_) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(currentaddr_19__FF_INPUT), .Q(currentaddr_19_) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(currentaddr_20__FF_INPUT), .Q(currentaddr_20_) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(currentaddr_21__FF_INPUT), .Q(currentaddr_21_) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(currentaddr_22__FF_INPUT), .Q(currentaddr_22_) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(currentaddr_23__FF_INPUT), .Q(currentaddr_23_) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(currentaddr_24__FF_INPUT), .Q(currentaddr_24_) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(currentaddr_25__FF_INPUT), .Q(currentaddr_25_) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(currentaddr_26__FF_INPUT), .Q(currentaddr_26_) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(currentaddr_27__FF_INPUT), .Q(currentaddr_27_) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(currentaddr_28__FF_INPUT), .Q(currentaddr_28_) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(currentaddr_29__FF_INPUT), .Q(currentaddr_29_) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(currentaddr_30__FF_INPUT), .Q(currentaddr_30_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(currentaddr_31__FF_INPUT), .Q(currentaddr_31_) );
	OR2X2 OR2X2_85 ( .A(addr[1]), .B(addr[0]), .Y(addr_decode__abc_3898_n21) );
	NAND2X1 NAND2X1_641 ( .A(addr[2]), .B(addr[3]), .Y(addr_decode__abc_3898_n22) );
	NOR2X1 NOR2X1_387 ( .A(addr_decode__abc_3898_n22), .B(addr_decode__abc_3898_n21), .Y(addr_ic) );
	INVX1 INVX1_115 ( .A(addr[0]), .Y(addr_decode__abc_3898_n24) );
	NAND2X1 NAND2X1_642 ( .A(addr[1]), .B(addr_decode__abc_3898_n24), .Y(addr_decode__abc_3898_n25) );
	NOR2X1 NOR2X1_388 ( .A(addr_decode__abc_3898_n22), .B(addr_decode__abc_3898_n25), .Y(addr_ia) );
	INVX1 INVX1_116 ( .A(addr[1]), .Y(addr_decode__abc_3898_n27_1) );
	NAND2X1 NAND2X1_643 ( .A(addr[0]), .B(addr_decode__abc_3898_n27_1), .Y(addr_decode__abc_3898_n28) );
	NOR2X1 NOR2X1_389 ( .A(addr_decode__abc_3898_n22), .B(addr_decode__abc_3898_n28), .Y(addr_ir) );
	NAND2X1 NAND2X1_644 ( .A(addr[1]), .B(addr[0]), .Y(addr_decode__abc_3898_n30) );
	NOR2X1 NOR2X1_390 ( .A(addr_decode__abc_3898_n22), .B(addr_decode__abc_3898_n30), .Y(addr_cr) );
	INVX1 INVX1_117 ( .A(addr[2]), .Y(addr_decode__abc_3898_n32) );
	NAND2X1 NAND2X1_645 ( .A(addr[3]), .B(addr_decode__abc_3898_n32), .Y(addr_decode__abc_3898_n33) );
	NOR2X1 NOR2X1_391 ( .A(addr_decode__abc_3898_n30), .B(addr_decode__abc_3898_n33), .Y(addr_sh) );
	INVX1 INVX1_118 ( .A(addr[3]), .Y(addr_decode__abc_3898_n35) );
	NAND2X1 NAND2X1_646 ( .A(addr[2]), .B(addr_decode__abc_3898_n35), .Y(addr_decode__abc_3898_n36) );
	NOR2X1 NOR2X1_392 ( .A(addr_decode__abc_3898_n21), .B(addr_decode__abc_3898_n36), .Y(addr_vb) );
	NOR2X1 NOR2X1_393 ( .A(addr_decode__abc_3898_n28), .B(addr_decode__abc_3898_n36), .Y(addr_vv) );
	OR2X2 OR2X2_86 ( .A(addr[2]), .B(addr[3]), .Y(addr_decode__abc_3898_n39_1) );
	NOR2X1 NOR2X1_394 ( .A(addr_decode__abc_3898_n39_1), .B(addr_decode__abc_3898_n28), .Y(addr_hv) );
	NOR2X1 NOR2X1_395 ( .A(addr_decode__abc_3898_n39_1), .B(addr_decode__abc_3898_n25), .Y(addr_hf) );
	NOR2X1 NOR2X1_396 ( .A(addr_decode__abc_3898_n21), .B(addr_decode__abc_3898_n33), .Y(addr_fl) );
	NOR2X1 NOR2X1_397 ( .A(addr_decode__abc_3898_n21), .B(addr_decode__abc_3898_n39_1), .Y(addr_hb) );
	NOR2X1 NOR2X1_398 ( .A(addr_decode__abc_3898_n30), .B(addr_decode__abc_3898_n36), .Y(addr_ve) );
	NOR2X1 NOR2X1_399 ( .A(addr_decode__abc_3898_n30), .B(addr_decode__abc_3898_n39_1), .Y(addr_he) );
	NOR2X1 NOR2X1_400 ( .A(addr_decode__abc_3898_n25), .B(addr_decode__abc_3898_n33), .Y(addr_sl) );
	NOR2X1 NOR2X1_401 ( .A(addr_decode__abc_3898_n28), .B(addr_decode__abc_3898_n33), .Y(addr_fh) );
	NOR2X1 NOR2X1_402 ( .A(addr_decode__abc_3898_n25), .B(addr_decode__abc_3898_n36), .Y(addr_vf) );
	INVX1 INVX1_119 ( .A(reg_cr_value_14_), .Y(reg_cr__abc_3798_n68_1) );
	INVX1 INVX1_120 ( .A(we), .Y(reg_cr__abc_3798_n69) );
	NAND2X1 NAND2X1_647 ( .A(addr_cr), .B(reg_cr__abc_3798_n69), .Y(reg_cr__abc_3798_n70_1) );
	NOR2X1 NOR2X1_403 ( .A(reg_cr__abc_3798_n68_1), .B(reg_cr__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_121 ( .A(reg_cr_value_13_), .Y(reg_cr__abc_3798_n72) );
	NOR2X1 NOR2X1_404 ( .A(reg_cr__abc_3798_n72), .B(reg_cr__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_122 ( .A(reg_cr_value_12_), .Y(reg_cr__abc_3798_n74_1) );
	NOR2X1 NOR2X1_405 ( .A(reg_cr__abc_3798_n74_1), .B(reg_cr__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_123 ( .A(reg_cr_value_11_), .Y(reg_cr__abc_3798_n76_1) );
	NOR2X1 NOR2X1_406 ( .A(reg_cr__abc_3798_n76_1), .B(reg_cr__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_124 ( .A(reg_cr_value_10_), .Y(reg_cr__abc_3798_n78) );
	NOR2X1 NOR2X1_407 ( .A(reg_cr__abc_3798_n78), .B(reg_cr__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_125 ( .A(reg_cr_value_9_), .Y(reg_cr__abc_3798_n80_1) );
	NOR2X1 NOR2X1_408 ( .A(reg_cr__abc_3798_n80_1), .B(reg_cr__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_126 ( .A(reg_cr_value_8_), .Y(reg_cr__abc_3798_n82_1) );
	NOR2X1 NOR2X1_409 ( .A(reg_cr__abc_3798_n82_1), .B(reg_cr__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_127 ( .A(reg_cr_value_7_), .Y(reg_cr__abc_3798_n84_1) );
	NOR2X1 NOR2X1_410 ( .A(reg_cr__abc_3798_n84_1), .B(reg_cr__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_128 ( .A(reg_cr_value_6_), .Y(reg_cr__abc_3798_n86) );
	NOR2X1 NOR2X1_411 ( .A(reg_cr__abc_3798_n86), .B(reg_cr__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_129 ( .A(reg_cr_value_5_), .Y(reg_cr__abc_3798_n88) );
	NOR2X1 NOR2X1_412 ( .A(reg_cr__abc_3798_n88), .B(reg_cr__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_130 ( .A(reg_cr_value_4_), .Y(reg_cr__abc_3798_n90) );
	NOR2X1 NOR2X1_413 ( .A(reg_cr__abc_3798_n90), .B(reg_cr__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_131 ( .A(reg_cr_value_3_), .Y(reg_cr__abc_3798_n92) );
	NOR2X1 NOR2X1_414 ( .A(reg_cr__abc_3798_n92), .B(reg_cr__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_132 ( .A(reg_cr_value_2_), .Y(reg_cr__abc_3798_n94) );
	NOR2X1 NOR2X1_415 ( .A(reg_cr__abc_3798_n94), .B(reg_cr__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_133 ( .A(reg_cr_value_1_), .Y(reg_cr__abc_3798_n96) );
	NOR2X1 NOR2X1_416 ( .A(reg_cr__abc_3798_n96), .B(reg_cr__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_134 ( .A(reg_cr_value_0_), .Y(reg_cr__abc_3798_n98) );
	NOR2X1 NOR2X1_417 ( .A(reg_cr__abc_3798_n98), .B(reg_cr__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_648 ( .A(we), .B(addr_cr), .Y(reg_cr__abc_3798_n100) );
	NOR2X1 NOR2X1_418 ( .A(reset), .B(reg_cr__abc_3798_n68_1), .Y(reg_cr__abc_3798_n101) );
	NAND2X1 NAND2X1_649 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n101), .Y(reg_cr__abc_3798_n102) );
	NAND2X1 NAND2X1_650 ( .A(gnd), .B(reset), .Y(reg_cr__abc_3798_n103) );
	NAND2X1 NAND2X1_651 ( .A(reg_cr__abc_3798_n103), .B(reg_cr__abc_3798_n102), .Y(reg_cr__abc_3798_n35) );
	NOR2X1 NOR2X1_419 ( .A(reset), .B(reg_cr__abc_3798_n72), .Y(reg_cr__abc_3798_n105) );
	NAND2X1 NAND2X1_652 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n105), .Y(reg_cr__abc_3798_n106) );
	NAND2X1 NAND2X1_653 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n107) );
	NAND2X1 NAND2X1_654 ( .A(reg_cr__abc_3798_n107), .B(reg_cr__abc_3798_n106), .Y(reg_cr__abc_3798_n38) );
	NOR2X1 NOR2X1_420 ( .A(reset), .B(reg_cr__abc_3798_n74_1), .Y(reg_cr__abc_3798_n109) );
	NAND2X1 NAND2X1_655 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n109), .Y(reg_cr__abc_3798_n110) );
	NAND2X1 NAND2X1_656 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n111) );
	NAND2X1 NAND2X1_657 ( .A(reg_cr__abc_3798_n111), .B(reg_cr__abc_3798_n110), .Y(reg_cr__abc_3798_n41) );
	NOR2X1 NOR2X1_421 ( .A(reset), .B(reg_cr__abc_3798_n76_1), .Y(reg_cr__abc_3798_n113) );
	NAND2X1 NAND2X1_658 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n113), .Y(reg_cr__abc_3798_n114) );
	NAND2X1 NAND2X1_659 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n115) );
	NAND2X1 NAND2X1_660 ( .A(reg_cr__abc_3798_n115), .B(reg_cr__abc_3798_n114), .Y(reg_cr__abc_3798_n44) );
	NOR2X1 NOR2X1_422 ( .A(reset), .B(reg_cr__abc_3798_n78), .Y(reg_cr__abc_3798_n117) );
	NAND2X1 NAND2X1_661 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n117), .Y(reg_cr__abc_3798_n118) );
	NAND2X1 NAND2X1_662 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n119) );
	NAND2X1 NAND2X1_663 ( .A(reg_cr__abc_3798_n119), .B(reg_cr__abc_3798_n118), .Y(reg_cr_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_423 ( .A(reset), .B(reg_cr__abc_3798_n80_1), .Y(reg_cr__abc_3798_n121) );
	NAND2X1 NAND2X1_664 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n121), .Y(reg_cr__abc_3798_n122) );
	NAND2X1 NAND2X1_665 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n123) );
	NAND2X1 NAND2X1_666 ( .A(reg_cr__abc_3798_n123), .B(reg_cr__abc_3798_n122), .Y(reg_cr_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_424 ( .A(reset), .B(reg_cr__abc_3798_n82_1), .Y(reg_cr__abc_3798_n125) );
	NAND2X1 NAND2X1_667 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n125), .Y(reg_cr__abc_3798_n126) );
	NAND2X1 NAND2X1_668 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n127) );
	NAND2X1 NAND2X1_669 ( .A(reg_cr__abc_3798_n127), .B(reg_cr__abc_3798_n126), .Y(reg_cr__abc_3798_n53) );
	NOR2X1 NOR2X1_425 ( .A(reset), .B(reg_cr__abc_3798_n84_1), .Y(reg_cr__abc_3798_n129) );
	NAND2X1 NAND2X1_670 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n129), .Y(reg_cr__abc_3798_n130) );
	NAND2X1 NAND2X1_671 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n131) );
	NAND2X1 NAND2X1_672 ( .A(reg_cr__abc_3798_n131), .B(reg_cr__abc_3798_n130), .Y(reg_cr__abc_3798_n56) );
	NOR2X1 NOR2X1_426 ( .A(reset), .B(reg_cr__abc_3798_n86), .Y(reg_cr__abc_3798_n133) );
	NAND2X1 NAND2X1_673 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n133), .Y(reg_cr__abc_3798_n134) );
	NAND2X1 NAND2X1_674 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n135) );
	NAND2X1 NAND2X1_675 ( .A(reg_cr__abc_3798_n135), .B(reg_cr__abc_3798_n134), .Y(reg_cr_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_427 ( .A(reset), .B(reg_cr__abc_3798_n88), .Y(reg_cr__abc_3798_n137) );
	NAND2X1 NAND2X1_676 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n137), .Y(reg_cr__abc_3798_n138) );
	NAND2X1 NAND2X1_677 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n139) );
	NAND2X1 NAND2X1_678 ( .A(reg_cr__abc_3798_n139), .B(reg_cr__abc_3798_n138), .Y(reg_cr_value_5__FF_INPUT) );
	NOR2X1 NOR2X1_428 ( .A(reset), .B(reg_cr__abc_3798_n90), .Y(reg_cr__abc_3798_n141) );
	NAND2X1 NAND2X1_679 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n141), .Y(reg_cr__abc_3798_n142) );
	NAND2X1 NAND2X1_680 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n143) );
	NAND2X1 NAND2X1_681 ( .A(reg_cr__abc_3798_n143), .B(reg_cr__abc_3798_n142), .Y(reg_cr_value_4__FF_INPUT) );
	NOR2X1 NOR2X1_429 ( .A(reset), .B(reg_cr__abc_3798_n92), .Y(reg_cr__abc_3798_n145) );
	NAND2X1 NAND2X1_682 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n145), .Y(reg_cr__abc_3798_n146) );
	NAND2X1 NAND2X1_683 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n147) );
	NAND2X1 NAND2X1_684 ( .A(reg_cr__abc_3798_n147), .B(reg_cr__abc_3798_n146), .Y(reg_cr_value_3__FF_INPUT) );
	NOR2X1 NOR2X1_430 ( .A(reset), .B(reg_cr__abc_3798_n94), .Y(reg_cr__abc_3798_n149) );
	NAND2X1 NAND2X1_685 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n149), .Y(reg_cr__abc_3798_n150) );
	NAND2X1 NAND2X1_686 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n151) );
	NAND2X1 NAND2X1_687 ( .A(reg_cr__abc_3798_n151), .B(reg_cr__abc_3798_n150), .Y(reg_cr_value_2__FF_INPUT) );
	NOR2X1 NOR2X1_431 ( .A(reset), .B(reg_cr__abc_3798_n96), .Y(reg_cr__abc_3798_n153) );
	NAND2X1 NAND2X1_688 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n153), .Y(reg_cr__abc_3798_n154) );
	NAND2X1 NAND2X1_689 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n155) );
	NAND2X1 NAND2X1_690 ( .A(reg_cr__abc_3798_n155), .B(reg_cr__abc_3798_n154), .Y(reg_cr_value_1__FF_INPUT) );
	NOR2X1 NOR2X1_432 ( .A(reset), .B(reg_cr__abc_3798_n98), .Y(reg_cr__abc_3798_n157) );
	NAND2X1 NAND2X1_691 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n157), .Y(reg_cr__abc_3798_n158) );
	NAND2X1 NAND2X1_692 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n159) );
	NAND2X1 NAND2X1_693 ( .A(reg_cr__abc_3798_n159), .B(reg_cr__abc_3798_n158), .Y(reg_cr_value_0__FF_INPUT) );
	INVX1 INVX1_135 ( .A(reg_cr_value_15_), .Y(reg_cr__abc_3798_n161) );
	NOR2X1 NOR2X1_433 ( .A(reset), .B(reg_cr__abc_3798_n161), .Y(reg_cr__abc_3798_n162) );
	NAND2X1 NAND2X1_694 ( .A(reg_cr__abc_3798_n100), .B(reg_cr__abc_3798_n162), .Y(reg_cr__abc_3798_n163) );
	NAND2X1 NAND2X1_695 ( .A(reset), .B(gnd), .Y(reg_cr__abc_3798_n164) );
	NAND2X1 NAND2X1_696 ( .A(reg_cr__abc_3798_n164), .B(reg_cr__abc_3798_n163), .Y(reg_cr_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_434 ( .A(reg_cr__abc_3798_n161), .B(reg_cr__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(reg_cr_value_0__FF_INPUT), .Q(reg_cr_value_0_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(reg_cr_value_1__FF_INPUT), .Q(reg_cr_value_1_) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(reg_cr_value_2__FF_INPUT), .Q(reg_cr_value_2_) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(reg_cr_value_3__FF_INPUT), .Q(reg_cr_value_3_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(reg_cr_value_4__FF_INPUT), .Q(reg_cr_value_4_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(reg_cr_value_5__FF_INPUT), .Q(reg_cr_value_5_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(reg_cr_value_6__FF_INPUT), .Q(reg_cr_value_6_) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(reg_cr__abc_3798_n56), .Q(reg_cr_value_7_) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(reg_cr__abc_3798_n53), .Q(reg_cr_value_8_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(reg_cr_value_9__FF_INPUT), .Q(reg_cr_value_9_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(reg_cr_value_10__FF_INPUT), .Q(reg_cr_value_10_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(reg_cr__abc_3798_n44), .Q(reg_cr_value_11_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(reg_cr__abc_3798_n41), .Q(reg_cr_value_12_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(reg_cr__abc_3798_n38), .Q(reg_cr_value_13_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(reg_cr__abc_3798_n35), .Q(reg_cr_value_14_) );
	DFFPOSX1 DFFPOSX1_81 ( .CLK(clk), .D(reg_cr_value_15__FF_INPUT), .Q(reg_cr_value_15_) );
	INVX1 INVX1_136 ( .A(reg_fh_value_14_), .Y(reg_fh__abc_3798_n68_1) );
	INVX1 INVX1_137 ( .A(we), .Y(reg_fh__abc_3798_n69) );
	NAND2X1 NAND2X1_697 ( .A(addr_fh), .B(reg_fh__abc_3798_n69), .Y(reg_fh__abc_3798_n70_1) );
	NOR2X1 NOR2X1_435 ( .A(reg_fh__abc_3798_n68_1), .B(reg_fh__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_138 ( .A(reg_fh_value_13_), .Y(reg_fh__abc_3798_n72) );
	NOR2X1 NOR2X1_436 ( .A(reg_fh__abc_3798_n72), .B(reg_fh__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_139 ( .A(reg_fh_value_12_), .Y(reg_fh__abc_3798_n74_1) );
	NOR2X1 NOR2X1_437 ( .A(reg_fh__abc_3798_n74_1), .B(reg_fh__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_140 ( .A(reg_fh_value_11_), .Y(reg_fh__abc_3798_n76_1) );
	NOR2X1 NOR2X1_438 ( .A(reg_fh__abc_3798_n76_1), .B(reg_fh__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_141 ( .A(reg_fh_value_10_), .Y(reg_fh__abc_3798_n78) );
	NOR2X1 NOR2X1_439 ( .A(reg_fh__abc_3798_n78), .B(reg_fh__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_142 ( .A(reg_fh_value_9_), .Y(reg_fh__abc_3798_n80_1) );
	NOR2X1 NOR2X1_440 ( .A(reg_fh__abc_3798_n80_1), .B(reg_fh__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_143 ( .A(reg_fh_value_8_), .Y(reg_fh__abc_3798_n82_1) );
	NOR2X1 NOR2X1_441 ( .A(reg_fh__abc_3798_n82_1), .B(reg_fh__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_144 ( .A(reg_fh_value_7_), .Y(reg_fh__abc_3798_n84_1) );
	NOR2X1 NOR2X1_442 ( .A(reg_fh__abc_3798_n84_1), .B(reg_fh__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_145 ( .A(reg_fh_value_6_), .Y(reg_fh__abc_3798_n86) );
	NOR2X1 NOR2X1_443 ( .A(reg_fh__abc_3798_n86), .B(reg_fh__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_146 ( .A(reg_fh_value_5_), .Y(reg_fh__abc_3798_n88) );
	NOR2X1 NOR2X1_444 ( .A(reg_fh__abc_3798_n88), .B(reg_fh__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_147 ( .A(reg_fh_value_4_), .Y(reg_fh__abc_3798_n90) );
	NOR2X1 NOR2X1_445 ( .A(reg_fh__abc_3798_n90), .B(reg_fh__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_148 ( .A(reg_fh_value_3_), .Y(reg_fh__abc_3798_n92) );
	NOR2X1 NOR2X1_446 ( .A(reg_fh__abc_3798_n92), .B(reg_fh__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_149 ( .A(reg_fh_value_2_), .Y(reg_fh__abc_3798_n94) );
	NOR2X1 NOR2X1_447 ( .A(reg_fh__abc_3798_n94), .B(reg_fh__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_150 ( .A(reg_fh_value_1_), .Y(reg_fh__abc_3798_n96) );
	NOR2X1 NOR2X1_448 ( .A(reg_fh__abc_3798_n96), .B(reg_fh__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_151 ( .A(reg_fh_value_0_), .Y(reg_fh__abc_3798_n98) );
	NOR2X1 NOR2X1_449 ( .A(reg_fh__abc_3798_n98), .B(reg_fh__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_698 ( .A(we), .B(addr_fh), .Y(reg_fh__abc_3798_n100) );
	NOR2X1 NOR2X1_450 ( .A(reset), .B(reg_fh__abc_3798_n68_1), .Y(reg_fh__abc_3798_n101) );
	NAND2X1 NAND2X1_699 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n101), .Y(reg_fh__abc_3798_n102) );
	NAND2X1 NAND2X1_700 ( .A(gnd), .B(reset), .Y(reg_fh__abc_3798_n103) );
	NAND2X1 NAND2X1_701 ( .A(reg_fh__abc_3798_n103), .B(reg_fh__abc_3798_n102), .Y(reg_fh__abc_3798_n35) );
	NOR2X1 NOR2X1_451 ( .A(reset), .B(reg_fh__abc_3798_n72), .Y(reg_fh__abc_3798_n105) );
	NAND2X1 NAND2X1_702 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n105), .Y(reg_fh__abc_3798_n106) );
	NAND2X1 NAND2X1_703 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n107) );
	NAND2X1 NAND2X1_704 ( .A(reg_fh__abc_3798_n107), .B(reg_fh__abc_3798_n106), .Y(reg_fh_value_13__FF_INPUT) );
	NOR2X1 NOR2X1_452 ( .A(reset), .B(reg_fh__abc_3798_n74_1), .Y(reg_fh__abc_3798_n109) );
	NAND2X1 NAND2X1_705 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n109), .Y(reg_fh__abc_3798_n110) );
	NAND2X1 NAND2X1_706 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n111) );
	NAND2X1 NAND2X1_707 ( .A(reg_fh__abc_3798_n111), .B(reg_fh__abc_3798_n110), .Y(reg_fh_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_453 ( .A(reset), .B(reg_fh__abc_3798_n76_1), .Y(reg_fh__abc_3798_n113) );
	NAND2X1 NAND2X1_708 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n113), .Y(reg_fh__abc_3798_n114) );
	NAND2X1 NAND2X1_709 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n115) );
	NAND2X1 NAND2X1_710 ( .A(reg_fh__abc_3798_n115), .B(reg_fh__abc_3798_n114), .Y(reg_fh__abc_3798_n44) );
	NOR2X1 NOR2X1_454 ( .A(reset), .B(reg_fh__abc_3798_n78), .Y(reg_fh__abc_3798_n117) );
	NAND2X1 NAND2X1_711 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n117), .Y(reg_fh__abc_3798_n118) );
	NAND2X1 NAND2X1_712 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n119) );
	NAND2X1 NAND2X1_713 ( .A(reg_fh__abc_3798_n119), .B(reg_fh__abc_3798_n118), .Y(reg_fh_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_455 ( .A(reset), .B(reg_fh__abc_3798_n80_1), .Y(reg_fh__abc_3798_n121) );
	NAND2X1 NAND2X1_714 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n121), .Y(reg_fh__abc_3798_n122) );
	NAND2X1 NAND2X1_715 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n123) );
	NAND2X1 NAND2X1_716 ( .A(reg_fh__abc_3798_n123), .B(reg_fh__abc_3798_n122), .Y(reg_fh_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_456 ( .A(reset), .B(reg_fh__abc_3798_n82_1), .Y(reg_fh__abc_3798_n125) );
	NAND2X1 NAND2X1_717 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n125), .Y(reg_fh__abc_3798_n126) );
	NAND2X1 NAND2X1_718 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n127) );
	NAND2X1 NAND2X1_719 ( .A(reg_fh__abc_3798_n127), .B(reg_fh__abc_3798_n126), .Y(reg_fh__abc_3798_n53) );
	NOR2X1 NOR2X1_457 ( .A(reset), .B(reg_fh__abc_3798_n84_1), .Y(reg_fh__abc_3798_n129) );
	NAND2X1 NAND2X1_720 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n129), .Y(reg_fh__abc_3798_n130) );
	NAND2X1 NAND2X1_721 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n131) );
	NAND2X1 NAND2X1_722 ( .A(reg_fh__abc_3798_n131), .B(reg_fh__abc_3798_n130), .Y(reg_fh_value_7__FF_INPUT) );
	NOR2X1 NOR2X1_458 ( .A(reset), .B(reg_fh__abc_3798_n86), .Y(reg_fh__abc_3798_n133) );
	NAND2X1 NAND2X1_723 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n133), .Y(reg_fh__abc_3798_n134) );
	NAND2X1 NAND2X1_724 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n135) );
	NAND2X1 NAND2X1_725 ( .A(reg_fh__abc_3798_n135), .B(reg_fh__abc_3798_n134), .Y(reg_fh_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_459 ( .A(reset), .B(reg_fh__abc_3798_n88), .Y(reg_fh__abc_3798_n137) );
	NAND2X1 NAND2X1_726 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n137), .Y(reg_fh__abc_3798_n138) );
	NAND2X1 NAND2X1_727 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n139) );
	NAND2X1 NAND2X1_728 ( .A(reg_fh__abc_3798_n139), .B(reg_fh__abc_3798_n138), .Y(reg_fh__abc_3798_n62) );
	NOR2X1 NOR2X1_460 ( .A(reset), .B(reg_fh__abc_3798_n90), .Y(reg_fh__abc_3798_n141) );
	NAND2X1 NAND2X1_729 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n141), .Y(reg_fh__abc_3798_n142) );
	NAND2X1 NAND2X1_730 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n143) );
	NAND2X1 NAND2X1_731 ( .A(reg_fh__abc_3798_n143), .B(reg_fh__abc_3798_n142), .Y(reg_fh_value_4__FF_INPUT) );
	NOR2X1 NOR2X1_461 ( .A(reset), .B(reg_fh__abc_3798_n92), .Y(reg_fh__abc_3798_n145) );
	NAND2X1 NAND2X1_732 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n145), .Y(reg_fh__abc_3798_n146) );
	NAND2X1 NAND2X1_733 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n147) );
	NAND2X1 NAND2X1_734 ( .A(reg_fh__abc_3798_n147), .B(reg_fh__abc_3798_n146), .Y(reg_fh__abc_3798_n68) );
	NOR2X1 NOR2X1_462 ( .A(reset), .B(reg_fh__abc_3798_n94), .Y(reg_fh__abc_3798_n149) );
	NAND2X1 NAND2X1_735 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n149), .Y(reg_fh__abc_3798_n150) );
	NAND2X1 NAND2X1_736 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n151) );
	NAND2X1 NAND2X1_737 ( .A(reg_fh__abc_3798_n151), .B(reg_fh__abc_3798_n150), .Y(reg_fh__abc_3798_n71) );
	NOR2X1 NOR2X1_463 ( .A(reset), .B(reg_fh__abc_3798_n96), .Y(reg_fh__abc_3798_n153) );
	NAND2X1 NAND2X1_738 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n153), .Y(reg_fh__abc_3798_n154) );
	NAND2X1 NAND2X1_739 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n155) );
	NAND2X1 NAND2X1_740 ( .A(reg_fh__abc_3798_n155), .B(reg_fh__abc_3798_n154), .Y(reg_fh__abc_3798_n74) );
	NOR2X1 NOR2X1_464 ( .A(reset), .B(reg_fh__abc_3798_n98), .Y(reg_fh__abc_3798_n157) );
	NAND2X1 NAND2X1_741 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n157), .Y(reg_fh__abc_3798_n158) );
	NAND2X1 NAND2X1_742 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n159) );
	NAND2X1 NAND2X1_743 ( .A(reg_fh__abc_3798_n159), .B(reg_fh__abc_3798_n158), .Y(reg_fh__abc_3798_n77) );
	INVX1 INVX1_152 ( .A(reg_fh_value_15_), .Y(reg_fh__abc_3798_n161) );
	NOR2X1 NOR2X1_465 ( .A(reset), .B(reg_fh__abc_3798_n161), .Y(reg_fh__abc_3798_n162) );
	NAND2X1 NAND2X1_744 ( .A(reg_fh__abc_3798_n100), .B(reg_fh__abc_3798_n162), .Y(reg_fh__abc_3798_n163) );
	NAND2X1 NAND2X1_745 ( .A(reset), .B(gnd), .Y(reg_fh__abc_3798_n164) );
	NAND2X1 NAND2X1_746 ( .A(reg_fh__abc_3798_n164), .B(reg_fh__abc_3798_n163), .Y(reg_fh_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_466 ( .A(reg_fh__abc_3798_n161), .B(reg_fh__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_82 ( .CLK(clk), .D(reg_fh__abc_3798_n77), .Q(reg_fh_value_0_) );
	DFFPOSX1 DFFPOSX1_83 ( .CLK(clk), .D(reg_fh__abc_3798_n74), .Q(reg_fh_value_1_) );
	DFFPOSX1 DFFPOSX1_84 ( .CLK(clk), .D(reg_fh__abc_3798_n71), .Q(reg_fh_value_2_) );
	DFFPOSX1 DFFPOSX1_85 ( .CLK(clk), .D(reg_fh__abc_3798_n68), .Q(reg_fh_value_3_) );
	DFFPOSX1 DFFPOSX1_86 ( .CLK(clk), .D(reg_fh_value_4__FF_INPUT), .Q(reg_fh_value_4_) );
	DFFPOSX1 DFFPOSX1_87 ( .CLK(clk), .D(reg_fh__abc_3798_n62), .Q(reg_fh_value_5_) );
	DFFPOSX1 DFFPOSX1_88 ( .CLK(clk), .D(reg_fh_value_6__FF_INPUT), .Q(reg_fh_value_6_) );
	DFFPOSX1 DFFPOSX1_89 ( .CLK(clk), .D(reg_fh_value_7__FF_INPUT), .Q(reg_fh_value_7_) );
	DFFPOSX1 DFFPOSX1_90 ( .CLK(clk), .D(reg_fh__abc_3798_n53), .Q(reg_fh_value_8_) );
	DFFPOSX1 DFFPOSX1_91 ( .CLK(clk), .D(reg_fh_value_9__FF_INPUT), .Q(reg_fh_value_9_) );
	DFFPOSX1 DFFPOSX1_92 ( .CLK(clk), .D(reg_fh_value_10__FF_INPUT), .Q(reg_fh_value_10_) );
	DFFPOSX1 DFFPOSX1_93 ( .CLK(clk), .D(reg_fh__abc_3798_n44), .Q(reg_fh_value_11_) );
	DFFPOSX1 DFFPOSX1_94 ( .CLK(clk), .D(reg_fh_value_12__FF_INPUT), .Q(reg_fh_value_12_) );
	DFFPOSX1 DFFPOSX1_95 ( .CLK(clk), .D(reg_fh_value_13__FF_INPUT), .Q(reg_fh_value_13_) );
	DFFPOSX1 DFFPOSX1_96 ( .CLK(clk), .D(reg_fh__abc_3798_n35), .Q(reg_fh_value_14_) );
	DFFPOSX1 DFFPOSX1_97 ( .CLK(clk), .D(reg_fh_value_15__FF_INPUT), .Q(reg_fh_value_15_) );
	INVX1 INVX1_153 ( .A(reg_fl_value_14_), .Y(reg_fl__abc_3798_n68_1) );
	INVX1 INVX1_154 ( .A(we), .Y(reg_fl__abc_3798_n69) );
	NAND2X1 NAND2X1_747 ( .A(addr_fl), .B(reg_fl__abc_3798_n69), .Y(reg_fl__abc_3798_n70_1) );
	NOR2X1 NOR2X1_467 ( .A(reg_fl__abc_3798_n68_1), .B(reg_fl__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_155 ( .A(reg_fl_value_13_), .Y(reg_fl__abc_3798_n72) );
	NOR2X1 NOR2X1_468 ( .A(reg_fl__abc_3798_n72), .B(reg_fl__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_156 ( .A(reg_fl_value_12_), .Y(reg_fl__abc_3798_n74_1) );
	NOR2X1 NOR2X1_469 ( .A(reg_fl__abc_3798_n74_1), .B(reg_fl__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_157 ( .A(reg_fl_value_11_), .Y(reg_fl__abc_3798_n76_1) );
	NOR2X1 NOR2X1_470 ( .A(reg_fl__abc_3798_n76_1), .B(reg_fl__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_158 ( .A(reg_fl_value_10_), .Y(reg_fl__abc_3798_n78) );
	NOR2X1 NOR2X1_471 ( .A(reg_fl__abc_3798_n78), .B(reg_fl__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_159 ( .A(reg_fl_value_9_), .Y(reg_fl__abc_3798_n80_1) );
	NOR2X1 NOR2X1_472 ( .A(reg_fl__abc_3798_n80_1), .B(reg_fl__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_160 ( .A(reg_fl_value_8_), .Y(reg_fl__abc_3798_n82_1) );
	NOR2X1 NOR2X1_473 ( .A(reg_fl__abc_3798_n82_1), .B(reg_fl__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_161 ( .A(reg_fl_value_7_), .Y(reg_fl__abc_3798_n84_1) );
	NOR2X1 NOR2X1_474 ( .A(reg_fl__abc_3798_n84_1), .B(reg_fl__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_162 ( .A(reg_fl_value_6_), .Y(reg_fl__abc_3798_n86) );
	NOR2X1 NOR2X1_475 ( .A(reg_fl__abc_3798_n86), .B(reg_fl__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_163 ( .A(reg_fl_value_5_), .Y(reg_fl__abc_3798_n88) );
	NOR2X1 NOR2X1_476 ( .A(reg_fl__abc_3798_n88), .B(reg_fl__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_164 ( .A(reg_fl_value_4_), .Y(reg_fl__abc_3798_n90) );
	NOR2X1 NOR2X1_477 ( .A(reg_fl__abc_3798_n90), .B(reg_fl__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_165 ( .A(reg_fl_value_3_), .Y(reg_fl__abc_3798_n92) );
	NOR2X1 NOR2X1_478 ( .A(reg_fl__abc_3798_n92), .B(reg_fl__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_166 ( .A(reg_fl_value_2_), .Y(reg_fl__abc_3798_n94) );
	NOR2X1 NOR2X1_479 ( .A(reg_fl__abc_3798_n94), .B(reg_fl__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_167 ( .A(reg_fl_value_1_), .Y(reg_fl__abc_3798_n96) );
	NOR2X1 NOR2X1_480 ( .A(reg_fl__abc_3798_n96), .B(reg_fl__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_168 ( .A(reg_fl_value_0_), .Y(reg_fl__abc_3798_n98) );
	NOR2X1 NOR2X1_481 ( .A(reg_fl__abc_3798_n98), .B(reg_fl__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_748 ( .A(we), .B(addr_fl), .Y(reg_fl__abc_3798_n100) );
	NOR2X1 NOR2X1_482 ( .A(reset), .B(reg_fl__abc_3798_n68_1), .Y(reg_fl__abc_3798_n101) );
	NAND2X1 NAND2X1_749 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n101), .Y(reg_fl__abc_3798_n102) );
	NAND2X1 NAND2X1_750 ( .A(gnd), .B(reset), .Y(reg_fl__abc_3798_n103) );
	NAND2X1 NAND2X1_751 ( .A(reg_fl__abc_3798_n103), .B(reg_fl__abc_3798_n102), .Y(reg_fl__abc_3798_n35) );
	NOR2X1 NOR2X1_483 ( .A(reset), .B(reg_fl__abc_3798_n72), .Y(reg_fl__abc_3798_n105) );
	NAND2X1 NAND2X1_752 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n105), .Y(reg_fl__abc_3798_n106) );
	NAND2X1 NAND2X1_753 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n107) );
	NAND2X1 NAND2X1_754 ( .A(reg_fl__abc_3798_n107), .B(reg_fl__abc_3798_n106), .Y(reg_fl__abc_3798_n38) );
	NOR2X1 NOR2X1_484 ( .A(reset), .B(reg_fl__abc_3798_n74_1), .Y(reg_fl__abc_3798_n109) );
	NAND2X1 NAND2X1_755 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n109), .Y(reg_fl__abc_3798_n110) );
	NAND2X1 NAND2X1_756 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n111) );
	NAND2X1 NAND2X1_757 ( .A(reg_fl__abc_3798_n111), .B(reg_fl__abc_3798_n110), .Y(reg_fl__abc_3798_n41) );
	NOR2X1 NOR2X1_485 ( .A(reset), .B(reg_fl__abc_3798_n76_1), .Y(reg_fl__abc_3798_n113) );
	NAND2X1 NAND2X1_758 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n113), .Y(reg_fl__abc_3798_n114) );
	NAND2X1 NAND2X1_759 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n115) );
	NAND2X1 NAND2X1_760 ( .A(reg_fl__abc_3798_n115), .B(reg_fl__abc_3798_n114), .Y(reg_fl__abc_3798_n44) );
	NOR2X1 NOR2X1_486 ( .A(reset), .B(reg_fl__abc_3798_n78), .Y(reg_fl__abc_3798_n117) );
	NAND2X1 NAND2X1_761 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n117), .Y(reg_fl__abc_3798_n118) );
	NAND2X1 NAND2X1_762 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n119) );
	NAND2X1 NAND2X1_763 ( .A(reg_fl__abc_3798_n119), .B(reg_fl__abc_3798_n118), .Y(reg_fl__abc_3798_n47) );
	NOR2X1 NOR2X1_487 ( .A(reset), .B(reg_fl__abc_3798_n80_1), .Y(reg_fl__abc_3798_n121) );
	NAND2X1 NAND2X1_764 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n121), .Y(reg_fl__abc_3798_n122) );
	NAND2X1 NAND2X1_765 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n123) );
	NAND2X1 NAND2X1_766 ( .A(reg_fl__abc_3798_n123), .B(reg_fl__abc_3798_n122), .Y(reg_fl__abc_3798_n50) );
	NOR2X1 NOR2X1_488 ( .A(reset), .B(reg_fl__abc_3798_n82_1), .Y(reg_fl__abc_3798_n125) );
	NAND2X1 NAND2X1_767 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n125), .Y(reg_fl__abc_3798_n126) );
	NAND2X1 NAND2X1_768 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n127) );
	NAND2X1 NAND2X1_769 ( .A(reg_fl__abc_3798_n127), .B(reg_fl__abc_3798_n126), .Y(reg_fl__abc_3798_n53) );
	NOR2X1 NOR2X1_489 ( .A(reset), .B(reg_fl__abc_3798_n84_1), .Y(reg_fl__abc_3798_n129) );
	NAND2X1 NAND2X1_770 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n129), .Y(reg_fl__abc_3798_n130) );
	NAND2X1 NAND2X1_771 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n131) );
	NAND2X1 NAND2X1_772 ( .A(reg_fl__abc_3798_n131), .B(reg_fl__abc_3798_n130), .Y(reg_fl__abc_3798_n56) );
	NOR2X1 NOR2X1_490 ( .A(reset), .B(reg_fl__abc_3798_n86), .Y(reg_fl__abc_3798_n133) );
	NAND2X1 NAND2X1_773 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n133), .Y(reg_fl__abc_3798_n134) );
	NAND2X1 NAND2X1_774 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n135) );
	NAND2X1 NAND2X1_775 ( .A(reg_fl__abc_3798_n135), .B(reg_fl__abc_3798_n134), .Y(reg_fl__abc_3798_n59) );
	NOR2X1 NOR2X1_491 ( .A(reset), .B(reg_fl__abc_3798_n88), .Y(reg_fl__abc_3798_n137) );
	NAND2X1 NAND2X1_776 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n137), .Y(reg_fl__abc_3798_n138) );
	NAND2X1 NAND2X1_777 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n139) );
	NAND2X1 NAND2X1_778 ( .A(reg_fl__abc_3798_n139), .B(reg_fl__abc_3798_n138), .Y(reg_fl__abc_3798_n62) );
	NOR2X1 NOR2X1_492 ( .A(reset), .B(reg_fl__abc_3798_n90), .Y(reg_fl__abc_3798_n141) );
	NAND2X1 NAND2X1_779 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n141), .Y(reg_fl__abc_3798_n142) );
	NAND2X1 NAND2X1_780 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n143) );
	NAND2X1 NAND2X1_781 ( .A(reg_fl__abc_3798_n143), .B(reg_fl__abc_3798_n142), .Y(reg_fl__abc_3798_n65) );
	NOR2X1 NOR2X1_493 ( .A(reset), .B(reg_fl__abc_3798_n92), .Y(reg_fl__abc_3798_n145) );
	NAND2X1 NAND2X1_782 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n145), .Y(reg_fl__abc_3798_n146) );
	NAND2X1 NAND2X1_783 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n147) );
	NAND2X1 NAND2X1_784 ( .A(reg_fl__abc_3798_n147), .B(reg_fl__abc_3798_n146), .Y(reg_fl__abc_3798_n68) );
	NOR2X1 NOR2X1_494 ( .A(reset), .B(reg_fl__abc_3798_n94), .Y(reg_fl__abc_3798_n149) );
	NAND2X1 NAND2X1_785 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n149), .Y(reg_fl__abc_3798_n150) );
	NAND2X1 NAND2X1_786 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n151) );
	NAND2X1 NAND2X1_787 ( .A(reg_fl__abc_3798_n151), .B(reg_fl__abc_3798_n150), .Y(reg_fl__abc_3798_n71) );
	NOR2X1 NOR2X1_495 ( .A(reset), .B(reg_fl__abc_3798_n96), .Y(reg_fl__abc_3798_n153) );
	NAND2X1 NAND2X1_788 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n153), .Y(reg_fl__abc_3798_n154) );
	NAND2X1 NAND2X1_789 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n155) );
	NAND2X1 NAND2X1_790 ( .A(reg_fl__abc_3798_n155), .B(reg_fl__abc_3798_n154), .Y(reg_fl__abc_3798_n74) );
	NOR2X1 NOR2X1_496 ( .A(reset), .B(reg_fl__abc_3798_n98), .Y(reg_fl__abc_3798_n157) );
	NAND2X1 NAND2X1_791 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n157), .Y(reg_fl__abc_3798_n158) );
	NAND2X1 NAND2X1_792 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n159) );
	NAND2X1 NAND2X1_793 ( .A(reg_fl__abc_3798_n159), .B(reg_fl__abc_3798_n158), .Y(reg_fl__abc_3798_n77) );
	INVX1 INVX1_169 ( .A(reg_fl_value_15_), .Y(reg_fl__abc_3798_n161) );
	NOR2X1 NOR2X1_497 ( .A(reset), .B(reg_fl__abc_3798_n161), .Y(reg_fl__abc_3798_n162) );
	NAND2X1 NAND2X1_794 ( .A(reg_fl__abc_3798_n100), .B(reg_fl__abc_3798_n162), .Y(reg_fl__abc_3798_n163) );
	NAND2X1 NAND2X1_795 ( .A(reset), .B(gnd), .Y(reg_fl__abc_3798_n164) );
	NAND2X1 NAND2X1_796 ( .A(reg_fl__abc_3798_n164), .B(reg_fl__abc_3798_n163), .Y(reg_fl__abc_3798_n81) );
	NOR2X1 NOR2X1_498 ( .A(reg_fl__abc_3798_n161), .B(reg_fl__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_98 ( .CLK(clk), .D(reg_fl__abc_3798_n77), .Q(reg_fl_value_0_) );
	DFFPOSX1 DFFPOSX1_99 ( .CLK(clk), .D(reg_fl__abc_3798_n74), .Q(reg_fl_value_1_) );
	DFFPOSX1 DFFPOSX1_100 ( .CLK(clk), .D(reg_fl__abc_3798_n71), .Q(reg_fl_value_2_) );
	DFFPOSX1 DFFPOSX1_101 ( .CLK(clk), .D(reg_fl__abc_3798_n68), .Q(reg_fl_value_3_) );
	DFFPOSX1 DFFPOSX1_102 ( .CLK(clk), .D(reg_fl__abc_3798_n65), .Q(reg_fl_value_4_) );
	DFFPOSX1 DFFPOSX1_103 ( .CLK(clk), .D(reg_fl__abc_3798_n62), .Q(reg_fl_value_5_) );
	DFFPOSX1 DFFPOSX1_104 ( .CLK(clk), .D(reg_fl__abc_3798_n59), .Q(reg_fl_value_6_) );
	DFFPOSX1 DFFPOSX1_105 ( .CLK(clk), .D(reg_fl__abc_3798_n56), .Q(reg_fl_value_7_) );
	DFFPOSX1 DFFPOSX1_106 ( .CLK(clk), .D(reg_fl__abc_3798_n53), .Q(reg_fl_value_8_) );
	DFFPOSX1 DFFPOSX1_107 ( .CLK(clk), .D(reg_fl__abc_3798_n50), .Q(reg_fl_value_9_) );
	DFFPOSX1 DFFPOSX1_108 ( .CLK(clk), .D(reg_fl__abc_3798_n47), .Q(reg_fl_value_10_) );
	DFFPOSX1 DFFPOSX1_109 ( .CLK(clk), .D(reg_fl__abc_3798_n44), .Q(reg_fl_value_11_) );
	DFFPOSX1 DFFPOSX1_110 ( .CLK(clk), .D(reg_fl__abc_3798_n41), .Q(reg_fl_value_12_) );
	DFFPOSX1 DFFPOSX1_111 ( .CLK(clk), .D(reg_fl__abc_3798_n38), .Q(reg_fl_value_13_) );
	DFFPOSX1 DFFPOSX1_112 ( .CLK(clk), .D(reg_fl__abc_3798_n35), .Q(reg_fl_value_14_) );
	DFFPOSX1 DFFPOSX1_113 ( .CLK(clk), .D(reg_fl__abc_3798_n81), .Q(reg_fl_value_15_) );
	INVX1 INVX1_170 ( .A(reg_hb_value_14_), .Y(reg_hb__abc_3798_n68_1) );
	INVX1 INVX1_171 ( .A(we), .Y(reg_hb__abc_3798_n69) );
	NAND2X1 NAND2X1_797 ( .A(addr_hb), .B(reg_hb__abc_3798_n69), .Y(reg_hb__abc_3798_n70_1) );
	NOR2X1 NOR2X1_499 ( .A(reg_hb__abc_3798_n68_1), .B(reg_hb__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_172 ( .A(reg_hb_value_13_), .Y(reg_hb__abc_3798_n72) );
	NOR2X1 NOR2X1_500 ( .A(reg_hb__abc_3798_n72), .B(reg_hb__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_173 ( .A(reg_hb_value_12_), .Y(reg_hb__abc_3798_n74_1) );
	NOR2X1 NOR2X1_501 ( .A(reg_hb__abc_3798_n74_1), .B(reg_hb__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_174 ( .A(reg_hb_value_11_), .Y(reg_hb__abc_3798_n76_1) );
	NOR2X1 NOR2X1_502 ( .A(reg_hb__abc_3798_n76_1), .B(reg_hb__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_175 ( .A(reg_hb_value_10_), .Y(reg_hb__abc_3798_n78) );
	NOR2X1 NOR2X1_503 ( .A(reg_hb__abc_3798_n78), .B(reg_hb__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_176 ( .A(reg_hb_value_9_), .Y(reg_hb__abc_3798_n80_1) );
	NOR2X1 NOR2X1_504 ( .A(reg_hb__abc_3798_n80_1), .B(reg_hb__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_177 ( .A(reg_hb_value_8_), .Y(reg_hb__abc_3798_n82_1) );
	NOR2X1 NOR2X1_505 ( .A(reg_hb__abc_3798_n82_1), .B(reg_hb__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_178 ( .A(reg_hb_value_7_), .Y(reg_hb__abc_3798_n84_1) );
	NOR2X1 NOR2X1_506 ( .A(reg_hb__abc_3798_n84_1), .B(reg_hb__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_179 ( .A(reg_hb_value_6_), .Y(reg_hb__abc_3798_n86) );
	NOR2X1 NOR2X1_507 ( .A(reg_hb__abc_3798_n86), .B(reg_hb__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_180 ( .A(reg_hb_value_5_), .Y(reg_hb__abc_3798_n88) );
	NOR2X1 NOR2X1_508 ( .A(reg_hb__abc_3798_n88), .B(reg_hb__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_181 ( .A(reg_hb_value_4_), .Y(reg_hb__abc_3798_n90) );
	NOR2X1 NOR2X1_509 ( .A(reg_hb__abc_3798_n90), .B(reg_hb__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_182 ( .A(reg_hb_value_3_), .Y(reg_hb__abc_3798_n92) );
	NOR2X1 NOR2X1_510 ( .A(reg_hb__abc_3798_n92), .B(reg_hb__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_183 ( .A(reg_hb_value_2_), .Y(reg_hb__abc_3798_n94) );
	NOR2X1 NOR2X1_511 ( .A(reg_hb__abc_3798_n94), .B(reg_hb__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_184 ( .A(reg_hb_value_1_), .Y(reg_hb__abc_3798_n96) );
	NOR2X1 NOR2X1_512 ( .A(reg_hb__abc_3798_n96), .B(reg_hb__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_185 ( .A(reg_hb_value_0_), .Y(reg_hb__abc_3798_n98) );
	NOR2X1 NOR2X1_513 ( .A(reg_hb__abc_3798_n98), .B(reg_hb__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_798 ( .A(we), .B(addr_hb), .Y(reg_hb__abc_3798_n100) );
	NOR2X1 NOR2X1_514 ( .A(reset), .B(reg_hb__abc_3798_n68_1), .Y(reg_hb__abc_3798_n101) );
	NAND2X1 NAND2X1_799 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n101), .Y(reg_hb__abc_3798_n102) );
	NAND2X1 NAND2X1_800 ( .A(gnd), .B(reset), .Y(reg_hb__abc_3798_n103) );
	NAND2X1 NAND2X1_801 ( .A(reg_hb__abc_3798_n103), .B(reg_hb__abc_3798_n102), .Y(reg_hb__abc_3798_n35) );
	NOR2X1 NOR2X1_515 ( .A(reset), .B(reg_hb__abc_3798_n72), .Y(reg_hb__abc_3798_n105) );
	NAND2X1 NAND2X1_802 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n105), .Y(reg_hb__abc_3798_n106) );
	NAND2X1 NAND2X1_803 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n107) );
	NAND2X1 NAND2X1_804 ( .A(reg_hb__abc_3798_n107), .B(reg_hb__abc_3798_n106), .Y(reg_hb__abc_3798_n38) );
	NOR2X1 NOR2X1_516 ( .A(reset), .B(reg_hb__abc_3798_n74_1), .Y(reg_hb__abc_3798_n109) );
	NAND2X1 NAND2X1_805 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n109), .Y(reg_hb__abc_3798_n110) );
	NAND2X1 NAND2X1_806 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n111) );
	NAND2X1 NAND2X1_807 ( .A(reg_hb__abc_3798_n111), .B(reg_hb__abc_3798_n110), .Y(reg_hb__abc_3798_n41) );
	NOR2X1 NOR2X1_517 ( .A(reset), .B(reg_hb__abc_3798_n76_1), .Y(reg_hb__abc_3798_n113) );
	NAND2X1 NAND2X1_808 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n113), .Y(reg_hb__abc_3798_n114) );
	NAND2X1 NAND2X1_809 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n115) );
	NAND2X1 NAND2X1_810 ( .A(reg_hb__abc_3798_n115), .B(reg_hb__abc_3798_n114), .Y(reg_hb__abc_3798_n44) );
	NOR2X1 NOR2X1_518 ( .A(reset), .B(reg_hb__abc_3798_n78), .Y(reg_hb__abc_3798_n117) );
	NAND2X1 NAND2X1_811 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n117), .Y(reg_hb__abc_3798_n118) );
	NAND2X1 NAND2X1_812 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n119) );
	NAND2X1 NAND2X1_813 ( .A(reg_hb__abc_3798_n119), .B(reg_hb__abc_3798_n118), .Y(reg_hb__abc_3798_n47) );
	NOR2X1 NOR2X1_519 ( .A(reset), .B(reg_hb__abc_3798_n80_1), .Y(reg_hb__abc_3798_n121) );
	NAND2X1 NAND2X1_814 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n121), .Y(reg_hb__abc_3798_n122) );
	NAND2X1 NAND2X1_815 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n123) );
	NAND2X1 NAND2X1_816 ( .A(reg_hb__abc_3798_n123), .B(reg_hb__abc_3798_n122), .Y(reg_hb__abc_3798_n50) );
	NOR2X1 NOR2X1_520 ( .A(reset), .B(reg_hb__abc_3798_n82_1), .Y(reg_hb__abc_3798_n125) );
	NAND2X1 NAND2X1_817 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n125), .Y(reg_hb__abc_3798_n126) );
	NAND2X1 NAND2X1_818 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n127) );
	NAND2X1 NAND2X1_819 ( .A(reg_hb__abc_3798_n127), .B(reg_hb__abc_3798_n126), .Y(reg_hb__abc_3798_n53) );
	NOR2X1 NOR2X1_521 ( .A(reset), .B(reg_hb__abc_3798_n84_1), .Y(reg_hb__abc_3798_n129) );
	NAND2X1 NAND2X1_820 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n129), .Y(reg_hb__abc_3798_n130) );
	NAND2X1 NAND2X1_821 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n131) );
	NAND2X1 NAND2X1_822 ( .A(reg_hb__abc_3798_n131), .B(reg_hb__abc_3798_n130), .Y(reg_hb__abc_3798_n56) );
	NOR2X1 NOR2X1_522 ( .A(reset), .B(reg_hb__abc_3798_n86), .Y(reg_hb__abc_3798_n133) );
	NAND2X1 NAND2X1_823 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n133), .Y(reg_hb__abc_3798_n134) );
	NAND2X1 NAND2X1_824 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n135) );
	NAND2X1 NAND2X1_825 ( .A(reg_hb__abc_3798_n135), .B(reg_hb__abc_3798_n134), .Y(reg_hb__abc_3798_n59) );
	NOR2X1 NOR2X1_523 ( .A(reset), .B(reg_hb__abc_3798_n88), .Y(reg_hb__abc_3798_n137) );
	NAND2X1 NAND2X1_826 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n137), .Y(reg_hb__abc_3798_n138) );
	NAND2X1 NAND2X1_827 ( .A(reset), .B(vdd), .Y(reg_hb__abc_3798_n139) );
	NAND2X1 NAND2X1_828 ( .A(reg_hb__abc_3798_n139), .B(reg_hb__abc_3798_n138), .Y(reg_hb__abc_3798_n62) );
	NOR2X1 NOR2X1_524 ( .A(reset), .B(reg_hb__abc_3798_n90), .Y(reg_hb__abc_3798_n141) );
	NAND2X1 NAND2X1_829 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n141), .Y(reg_hb__abc_3798_n142) );
	NAND2X1 NAND2X1_830 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n143) );
	NAND2X1 NAND2X1_831 ( .A(reg_hb__abc_3798_n143), .B(reg_hb__abc_3798_n142), .Y(reg_hb__abc_3798_n65) );
	NOR2X1 NOR2X1_525 ( .A(reset), .B(reg_hb__abc_3798_n92), .Y(reg_hb__abc_3798_n145) );
	NAND2X1 NAND2X1_832 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n145), .Y(reg_hb__abc_3798_n146) );
	NAND2X1 NAND2X1_833 ( .A(reset), .B(vdd), .Y(reg_hb__abc_3798_n147) );
	NAND2X1 NAND2X1_834 ( .A(reg_hb__abc_3798_n147), .B(reg_hb__abc_3798_n146), .Y(reg_hb__abc_3798_n68) );
	NOR2X1 NOR2X1_526 ( .A(reset), .B(reg_hb__abc_3798_n94), .Y(reg_hb__abc_3798_n149) );
	NAND2X1 NAND2X1_835 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n149), .Y(reg_hb__abc_3798_n150) );
	NAND2X1 NAND2X1_836 ( .A(reset), .B(vdd), .Y(reg_hb__abc_3798_n151) );
	NAND2X1 NAND2X1_837 ( .A(reg_hb__abc_3798_n151), .B(reg_hb__abc_3798_n150), .Y(reg_hb__abc_3798_n71) );
	NOR2X1 NOR2X1_527 ( .A(reset), .B(reg_hb__abc_3798_n96), .Y(reg_hb__abc_3798_n153) );
	NAND2X1 NAND2X1_838 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n153), .Y(reg_hb__abc_3798_n154) );
	NAND2X1 NAND2X1_839 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n155) );
	NAND2X1 NAND2X1_840 ( .A(reg_hb__abc_3798_n155), .B(reg_hb__abc_3798_n154), .Y(reg_hb__abc_3798_n74) );
	NOR2X1 NOR2X1_528 ( .A(reset), .B(reg_hb__abc_3798_n98), .Y(reg_hb__abc_3798_n157) );
	NAND2X1 NAND2X1_841 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n157), .Y(reg_hb__abc_3798_n158) );
	NAND2X1 NAND2X1_842 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n159) );
	NAND2X1 NAND2X1_843 ( .A(reg_hb__abc_3798_n159), .B(reg_hb__abc_3798_n158), .Y(reg_hb__abc_3798_n77) );
	INVX1 INVX1_186 ( .A(reg_hb_value_15_), .Y(reg_hb__abc_3798_n161) );
	NOR2X1 NOR2X1_529 ( .A(reset), .B(reg_hb__abc_3798_n161), .Y(reg_hb__abc_3798_n162) );
	NAND2X1 NAND2X1_844 ( .A(reg_hb__abc_3798_n100), .B(reg_hb__abc_3798_n162), .Y(reg_hb__abc_3798_n163) );
	NAND2X1 NAND2X1_845 ( .A(reset), .B(gnd), .Y(reg_hb__abc_3798_n164) );
	NAND2X1 NAND2X1_846 ( .A(reg_hb__abc_3798_n164), .B(reg_hb__abc_3798_n163), .Y(reg_hb__abc_3798_n81) );
	NOR2X1 NOR2X1_530 ( .A(reg_hb__abc_3798_n161), .B(reg_hb__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_114 ( .CLK(clk), .D(reg_hb__abc_3798_n77), .Q(reg_hb_value_0_) );
	DFFPOSX1 DFFPOSX1_115 ( .CLK(clk), .D(reg_hb__abc_3798_n74), .Q(reg_hb_value_1_) );
	DFFPOSX1 DFFPOSX1_116 ( .CLK(clk), .D(reg_hb__abc_3798_n71), .Q(reg_hb_value_2_) );
	DFFPOSX1 DFFPOSX1_117 ( .CLK(clk), .D(reg_hb__abc_3798_n68), .Q(reg_hb_value_3_) );
	DFFPOSX1 DFFPOSX1_118 ( .CLK(clk), .D(reg_hb__abc_3798_n65), .Q(reg_hb_value_4_) );
	DFFPOSX1 DFFPOSX1_119 ( .CLK(clk), .D(reg_hb__abc_3798_n62), .Q(reg_hb_value_5_) );
	DFFPOSX1 DFFPOSX1_120 ( .CLK(clk), .D(reg_hb__abc_3798_n59), .Q(reg_hb_value_6_) );
	DFFPOSX1 DFFPOSX1_121 ( .CLK(clk), .D(reg_hb__abc_3798_n56), .Q(reg_hb_value_7_) );
	DFFPOSX1 DFFPOSX1_122 ( .CLK(clk), .D(reg_hb__abc_3798_n53), .Q(reg_hb_value_8_) );
	DFFPOSX1 DFFPOSX1_123 ( .CLK(clk), .D(reg_hb__abc_3798_n50), .Q(reg_hb_value_9_) );
	DFFPOSX1 DFFPOSX1_124 ( .CLK(clk), .D(reg_hb__abc_3798_n47), .Q(reg_hb_value_10_) );
	DFFPOSX1 DFFPOSX1_125 ( .CLK(clk), .D(reg_hb__abc_3798_n44), .Q(reg_hb_value_11_) );
	DFFPOSX1 DFFPOSX1_126 ( .CLK(clk), .D(reg_hb__abc_3798_n41), .Q(reg_hb_value_12_) );
	DFFPOSX1 DFFPOSX1_127 ( .CLK(clk), .D(reg_hb__abc_3798_n38), .Q(reg_hb_value_13_) );
	DFFPOSX1 DFFPOSX1_128 ( .CLK(clk), .D(reg_hb__abc_3798_n35), .Q(reg_hb_value_14_) );
	DFFPOSX1 DFFPOSX1_129 ( .CLK(clk), .D(reg_hb__abc_3798_n81), .Q(reg_hb_value_15_) );
	INVX1 INVX1_187 ( .A(reg_he_value_14_), .Y(reg_he__abc_3798_n68_1) );
	INVX1 INVX1_188 ( .A(we), .Y(reg_he__abc_3798_n69) );
	NAND2X1 NAND2X1_847 ( .A(addr_he), .B(reg_he__abc_3798_n69), .Y(reg_he__abc_3798_n70_1) );
	NOR2X1 NOR2X1_531 ( .A(reg_he__abc_3798_n68_1), .B(reg_he__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_189 ( .A(reg_he_value_13_), .Y(reg_he__abc_3798_n72) );
	NOR2X1 NOR2X1_532 ( .A(reg_he__abc_3798_n72), .B(reg_he__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_190 ( .A(reg_he_value_12_), .Y(reg_he__abc_3798_n74_1) );
	NOR2X1 NOR2X1_533 ( .A(reg_he__abc_3798_n74_1), .B(reg_he__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_191 ( .A(reg_he_value_11_), .Y(reg_he__abc_3798_n76_1) );
	NOR2X1 NOR2X1_534 ( .A(reg_he__abc_3798_n76_1), .B(reg_he__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_192 ( .A(reg_he_value_10_), .Y(reg_he__abc_3798_n78) );
	NOR2X1 NOR2X1_535 ( .A(reg_he__abc_3798_n78), .B(reg_he__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_193 ( .A(reg_he_value_9_), .Y(reg_he__abc_3798_n80_1) );
	NOR2X1 NOR2X1_536 ( .A(reg_he__abc_3798_n80_1), .B(reg_he__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_194 ( .A(reg_he_value_8_), .Y(reg_he__abc_3798_n82_1) );
	NOR2X1 NOR2X1_537 ( .A(reg_he__abc_3798_n82_1), .B(reg_he__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_195 ( .A(reg_he_value_7_), .Y(reg_he__abc_3798_n84_1) );
	NOR2X1 NOR2X1_538 ( .A(reg_he__abc_3798_n84_1), .B(reg_he__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_196 ( .A(reg_he_value_6_), .Y(reg_he__abc_3798_n86) );
	NOR2X1 NOR2X1_539 ( .A(reg_he__abc_3798_n86), .B(reg_he__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_197 ( .A(reg_he_value_5_), .Y(reg_he__abc_3798_n88) );
	NOR2X1 NOR2X1_540 ( .A(reg_he__abc_3798_n88), .B(reg_he__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_198 ( .A(reg_he_value_4_), .Y(reg_he__abc_3798_n90) );
	NOR2X1 NOR2X1_541 ( .A(reg_he__abc_3798_n90), .B(reg_he__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_199 ( .A(reg_he_value_3_), .Y(reg_he__abc_3798_n92) );
	NOR2X1 NOR2X1_542 ( .A(reg_he__abc_3798_n92), .B(reg_he__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_200 ( .A(reg_he_value_2_), .Y(reg_he__abc_3798_n94) );
	NOR2X1 NOR2X1_543 ( .A(reg_he__abc_3798_n94), .B(reg_he__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_201 ( .A(reg_he_value_1_), .Y(reg_he__abc_3798_n96) );
	NOR2X1 NOR2X1_544 ( .A(reg_he__abc_3798_n96), .B(reg_he__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_202 ( .A(reg_he_value_0_), .Y(reg_he__abc_3798_n98) );
	NOR2X1 NOR2X1_545 ( .A(reg_he__abc_3798_n98), .B(reg_he__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_848 ( .A(we), .B(addr_he), .Y(reg_he__abc_3798_n100) );
	NOR2X1 NOR2X1_546 ( .A(reset), .B(reg_he__abc_3798_n68_1), .Y(reg_he__abc_3798_n101) );
	NAND2X1 NAND2X1_849 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n101), .Y(reg_he__abc_3798_n102) );
	NAND2X1 NAND2X1_850 ( .A(gnd), .B(reset), .Y(reg_he__abc_3798_n103) );
	NAND2X1 NAND2X1_851 ( .A(reg_he__abc_3798_n103), .B(reg_he__abc_3798_n102), .Y(reg_he_value_14__FF_INPUT) );
	NOR2X1 NOR2X1_547 ( .A(reset), .B(reg_he__abc_3798_n72), .Y(reg_he__abc_3798_n105) );
	NAND2X1 NAND2X1_852 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n105), .Y(reg_he__abc_3798_n106) );
	NAND2X1 NAND2X1_853 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n107) );
	NAND2X1 NAND2X1_854 ( .A(reg_he__abc_3798_n107), .B(reg_he__abc_3798_n106), .Y(reg_he__abc_3798_n38) );
	NOR2X1 NOR2X1_548 ( .A(reset), .B(reg_he__abc_3798_n74_1), .Y(reg_he__abc_3798_n109) );
	NAND2X1 NAND2X1_855 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n109), .Y(reg_he__abc_3798_n110) );
	NAND2X1 NAND2X1_856 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n111) );
	NAND2X1 NAND2X1_857 ( .A(reg_he__abc_3798_n111), .B(reg_he__abc_3798_n110), .Y(reg_he_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_549 ( .A(reset), .B(reg_he__abc_3798_n76_1), .Y(reg_he__abc_3798_n113) );
	NAND2X1 NAND2X1_858 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n113), .Y(reg_he__abc_3798_n114) );
	NAND2X1 NAND2X1_859 ( .A(reset), .B(vdd), .Y(reg_he__abc_3798_n115) );
	NAND2X1 NAND2X1_860 ( .A(reg_he__abc_3798_n115), .B(reg_he__abc_3798_n114), .Y(reg_he_value_11__FF_INPUT) );
	NOR2X1 NOR2X1_550 ( .A(reset), .B(reg_he__abc_3798_n78), .Y(reg_he__abc_3798_n117) );
	NAND2X1 NAND2X1_861 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n117), .Y(reg_he__abc_3798_n118) );
	NAND2X1 NAND2X1_862 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n119) );
	NAND2X1 NAND2X1_863 ( .A(reg_he__abc_3798_n119), .B(reg_he__abc_3798_n118), .Y(reg_he_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_551 ( .A(reset), .B(reg_he__abc_3798_n80_1), .Y(reg_he__abc_3798_n121) );
	NAND2X1 NAND2X1_864 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n121), .Y(reg_he__abc_3798_n122) );
	NAND2X1 NAND2X1_865 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n123) );
	NAND2X1 NAND2X1_866 ( .A(reg_he__abc_3798_n123), .B(reg_he__abc_3798_n122), .Y(reg_he__abc_3798_n50) );
	NOR2X1 NOR2X1_552 ( .A(reset), .B(reg_he__abc_3798_n82_1), .Y(reg_he__abc_3798_n125) );
	NAND2X1 NAND2X1_867 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n125), .Y(reg_he__abc_3798_n126) );
	NAND2X1 NAND2X1_868 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n127) );
	NAND2X1 NAND2X1_869 ( .A(reg_he__abc_3798_n127), .B(reg_he__abc_3798_n126), .Y(reg_he__abc_3798_n53) );
	NOR2X1 NOR2X1_553 ( .A(reset), .B(reg_he__abc_3798_n84_1), .Y(reg_he__abc_3798_n129) );
	NAND2X1 NAND2X1_870 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n129), .Y(reg_he__abc_3798_n130) );
	NAND2X1 NAND2X1_871 ( .A(reset), .B(vdd), .Y(reg_he__abc_3798_n131) );
	NAND2X1 NAND2X1_872 ( .A(reg_he__abc_3798_n131), .B(reg_he__abc_3798_n130), .Y(reg_he__abc_3798_n56) );
	NOR2X1 NOR2X1_554 ( .A(reset), .B(reg_he__abc_3798_n86), .Y(reg_he__abc_3798_n133) );
	NAND2X1 NAND2X1_873 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n133), .Y(reg_he__abc_3798_n134) );
	NAND2X1 NAND2X1_874 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n135) );
	NAND2X1 NAND2X1_875 ( .A(reg_he__abc_3798_n135), .B(reg_he__abc_3798_n134), .Y(reg_he__abc_3798_n59) );
	NOR2X1 NOR2X1_555 ( .A(reset), .B(reg_he__abc_3798_n88), .Y(reg_he__abc_3798_n137) );
	NAND2X1 NAND2X1_876 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n137), .Y(reg_he__abc_3798_n138) );
	NAND2X1 NAND2X1_877 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n139) );
	NAND2X1 NAND2X1_878 ( .A(reg_he__abc_3798_n139), .B(reg_he__abc_3798_n138), .Y(reg_he__abc_3798_n62) );
	NOR2X1 NOR2X1_556 ( .A(reset), .B(reg_he__abc_3798_n90), .Y(reg_he__abc_3798_n141) );
	NAND2X1 NAND2X1_879 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n141), .Y(reg_he__abc_3798_n142) );
	NAND2X1 NAND2X1_880 ( .A(reset), .B(vdd), .Y(reg_he__abc_3798_n143) );
	NAND2X1 NAND2X1_881 ( .A(reg_he__abc_3798_n143), .B(reg_he__abc_3798_n142), .Y(reg_he__abc_3798_n65) );
	NOR2X1 NOR2X1_557 ( .A(reset), .B(reg_he__abc_3798_n92), .Y(reg_he__abc_3798_n145) );
	NAND2X1 NAND2X1_882 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n145), .Y(reg_he__abc_3798_n146) );
	NAND2X1 NAND2X1_883 ( .A(reset), .B(vdd), .Y(reg_he__abc_3798_n147) );
	NAND2X1 NAND2X1_884 ( .A(reg_he__abc_3798_n147), .B(reg_he__abc_3798_n146), .Y(reg_he__abc_3798_n68) );
	NOR2X1 NOR2X1_558 ( .A(reset), .B(reg_he__abc_3798_n94), .Y(reg_he__abc_3798_n149) );
	NAND2X1 NAND2X1_885 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n149), .Y(reg_he__abc_3798_n150) );
	NAND2X1 NAND2X1_886 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n151) );
	NAND2X1 NAND2X1_887 ( .A(reg_he__abc_3798_n151), .B(reg_he__abc_3798_n150), .Y(reg_he__abc_3798_n71) );
	NOR2X1 NOR2X1_559 ( .A(reset), .B(reg_he__abc_3798_n96), .Y(reg_he__abc_3798_n153) );
	NAND2X1 NAND2X1_888 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n153), .Y(reg_he__abc_3798_n154) );
	NAND2X1 NAND2X1_889 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n155) );
	NAND2X1 NAND2X1_890 ( .A(reg_he__abc_3798_n155), .B(reg_he__abc_3798_n154), .Y(reg_he_value_1__FF_INPUT) );
	NOR2X1 NOR2X1_560 ( .A(reset), .B(reg_he__abc_3798_n98), .Y(reg_he__abc_3798_n157) );
	NAND2X1 NAND2X1_891 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n157), .Y(reg_he__abc_3798_n158) );
	NAND2X1 NAND2X1_892 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n159) );
	NAND2X1 NAND2X1_893 ( .A(reg_he__abc_3798_n159), .B(reg_he__abc_3798_n158), .Y(reg_he_value_0__FF_INPUT) );
	INVX1 INVX1_203 ( .A(reg_he_value_15_), .Y(reg_he__abc_3798_n161) );
	NOR2X1 NOR2X1_561 ( .A(reset), .B(reg_he__abc_3798_n161), .Y(reg_he__abc_3798_n162) );
	NAND2X1 NAND2X1_894 ( .A(reg_he__abc_3798_n100), .B(reg_he__abc_3798_n162), .Y(reg_he__abc_3798_n163) );
	NAND2X1 NAND2X1_895 ( .A(reset), .B(gnd), .Y(reg_he__abc_3798_n164) );
	NAND2X1 NAND2X1_896 ( .A(reg_he__abc_3798_n164), .B(reg_he__abc_3798_n163), .Y(reg_he_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_562 ( .A(reg_he__abc_3798_n161), .B(reg_he__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_130 ( .CLK(clk), .D(reg_he_value_0__FF_INPUT), .Q(reg_he_value_0_) );
	DFFPOSX1 DFFPOSX1_131 ( .CLK(clk), .D(reg_he_value_1__FF_INPUT), .Q(reg_he_value_1_) );
	DFFPOSX1 DFFPOSX1_132 ( .CLK(clk), .D(reg_he__abc_3798_n71), .Q(reg_he_value_2_) );
	DFFPOSX1 DFFPOSX1_133 ( .CLK(clk), .D(reg_he__abc_3798_n68), .Q(reg_he_value_3_) );
	DFFPOSX1 DFFPOSX1_134 ( .CLK(clk), .D(reg_he__abc_3798_n65), .Q(reg_he_value_4_) );
	DFFPOSX1 DFFPOSX1_135 ( .CLK(clk), .D(reg_he__abc_3798_n62), .Q(reg_he_value_5_) );
	DFFPOSX1 DFFPOSX1_136 ( .CLK(clk), .D(reg_he__abc_3798_n59), .Q(reg_he_value_6_) );
	DFFPOSX1 DFFPOSX1_137 ( .CLK(clk), .D(reg_he__abc_3798_n56), .Q(reg_he_value_7_) );
	DFFPOSX1 DFFPOSX1_138 ( .CLK(clk), .D(reg_he__abc_3798_n53), .Q(reg_he_value_8_) );
	DFFPOSX1 DFFPOSX1_139 ( .CLK(clk), .D(reg_he__abc_3798_n50), .Q(reg_he_value_9_) );
	DFFPOSX1 DFFPOSX1_140 ( .CLK(clk), .D(reg_he_value_10__FF_INPUT), .Q(reg_he_value_10_) );
	DFFPOSX1 DFFPOSX1_141 ( .CLK(clk), .D(reg_he_value_11__FF_INPUT), .Q(reg_he_value_11_) );
	DFFPOSX1 DFFPOSX1_142 ( .CLK(clk), .D(reg_he_value_12__FF_INPUT), .Q(reg_he_value_12_) );
	DFFPOSX1 DFFPOSX1_143 ( .CLK(clk), .D(reg_he__abc_3798_n38), .Q(reg_he_value_13_) );
	DFFPOSX1 DFFPOSX1_144 ( .CLK(clk), .D(reg_he_value_14__FF_INPUT), .Q(reg_he_value_14_) );
	DFFPOSX1 DFFPOSX1_145 ( .CLK(clk), .D(reg_he_value_15__FF_INPUT), .Q(reg_he_value_15_) );
	INVX1 INVX1_204 ( .A(reg_hf_value_14_), .Y(reg_hf__abc_3798_n68_1) );
	INVX1 INVX1_205 ( .A(we), .Y(reg_hf__abc_3798_n69) );
	NAND2X1 NAND2X1_897 ( .A(addr_hf), .B(reg_hf__abc_3798_n69), .Y(reg_hf__abc_3798_n70_1) );
	NOR2X1 NOR2X1_563 ( .A(reg_hf__abc_3798_n68_1), .B(reg_hf__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_206 ( .A(reg_hf_value_13_), .Y(reg_hf__abc_3798_n72) );
	NOR2X1 NOR2X1_564 ( .A(reg_hf__abc_3798_n72), .B(reg_hf__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_207 ( .A(reg_hf_value_12_), .Y(reg_hf__abc_3798_n74_1) );
	NOR2X1 NOR2X1_565 ( .A(reg_hf__abc_3798_n74_1), .B(reg_hf__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_208 ( .A(reg_hf_value_11_), .Y(reg_hf__abc_3798_n76_1) );
	NOR2X1 NOR2X1_566 ( .A(reg_hf__abc_3798_n76_1), .B(reg_hf__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_209 ( .A(reg_hf_value_10_), .Y(reg_hf__abc_3798_n78) );
	NOR2X1 NOR2X1_567 ( .A(reg_hf__abc_3798_n78), .B(reg_hf__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_210 ( .A(reg_hf_value_9_), .Y(reg_hf__abc_3798_n80_1) );
	NOR2X1 NOR2X1_568 ( .A(reg_hf__abc_3798_n80_1), .B(reg_hf__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_211 ( .A(reg_hf_value_8_), .Y(reg_hf__abc_3798_n82_1) );
	NOR2X1 NOR2X1_569 ( .A(reg_hf__abc_3798_n82_1), .B(reg_hf__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_212 ( .A(reg_hf_value_7_), .Y(reg_hf__abc_3798_n84_1) );
	NOR2X1 NOR2X1_570 ( .A(reg_hf__abc_3798_n84_1), .B(reg_hf__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_213 ( .A(reg_hf_value_6_), .Y(reg_hf__abc_3798_n86) );
	NOR2X1 NOR2X1_571 ( .A(reg_hf__abc_3798_n86), .B(reg_hf__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_214 ( .A(reg_hf_value_5_), .Y(reg_hf__abc_3798_n88) );
	NOR2X1 NOR2X1_572 ( .A(reg_hf__abc_3798_n88), .B(reg_hf__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_215 ( .A(reg_hf_value_4_), .Y(reg_hf__abc_3798_n90) );
	NOR2X1 NOR2X1_573 ( .A(reg_hf__abc_3798_n90), .B(reg_hf__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_216 ( .A(reg_hf_value_3_), .Y(reg_hf__abc_3798_n92) );
	NOR2X1 NOR2X1_574 ( .A(reg_hf__abc_3798_n92), .B(reg_hf__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_217 ( .A(reg_hf_value_2_), .Y(reg_hf__abc_3798_n94) );
	NOR2X1 NOR2X1_575 ( .A(reg_hf__abc_3798_n94), .B(reg_hf__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_218 ( .A(reg_hf_value_1_), .Y(reg_hf__abc_3798_n96) );
	NOR2X1 NOR2X1_576 ( .A(reg_hf__abc_3798_n96), .B(reg_hf__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_219 ( .A(reg_hf_value_0_), .Y(reg_hf__abc_3798_n98) );
	NOR2X1 NOR2X1_577 ( .A(reg_hf__abc_3798_n98), .B(reg_hf__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_898 ( .A(we), .B(addr_hf), .Y(reg_hf__abc_3798_n100) );
	NOR2X1 NOR2X1_578 ( .A(reset), .B(reg_hf__abc_3798_n68_1), .Y(reg_hf__abc_3798_n101) );
	NAND2X1 NAND2X1_899 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n101), .Y(reg_hf__abc_3798_n102) );
	NAND2X1 NAND2X1_900 ( .A(gnd), .B(reset), .Y(reg_hf__abc_3798_n103) );
	NAND2X1 NAND2X1_901 ( .A(reg_hf__abc_3798_n103), .B(reg_hf__abc_3798_n102), .Y(reg_hf_value_14__FF_INPUT) );
	NOR2X1 NOR2X1_579 ( .A(reset), .B(reg_hf__abc_3798_n72), .Y(reg_hf__abc_3798_n105) );
	NAND2X1 NAND2X1_902 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n105), .Y(reg_hf__abc_3798_n106) );
	NAND2X1 NAND2X1_903 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n107) );
	NAND2X1 NAND2X1_904 ( .A(reg_hf__abc_3798_n107), .B(reg_hf__abc_3798_n106), .Y(reg_hf_value_13__FF_INPUT) );
	NOR2X1 NOR2X1_580 ( .A(reset), .B(reg_hf__abc_3798_n74_1), .Y(reg_hf__abc_3798_n109) );
	NAND2X1 NAND2X1_905 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n109), .Y(reg_hf__abc_3798_n110) );
	NAND2X1 NAND2X1_906 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n111) );
	NAND2X1 NAND2X1_907 ( .A(reg_hf__abc_3798_n111), .B(reg_hf__abc_3798_n110), .Y(reg_hf_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_581 ( .A(reset), .B(reg_hf__abc_3798_n76_1), .Y(reg_hf__abc_3798_n113) );
	NAND2X1 NAND2X1_908 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n113), .Y(reg_hf__abc_3798_n114) );
	NAND2X1 NAND2X1_909 ( .A(reset), .B(vdd), .Y(reg_hf__abc_3798_n115) );
	NAND2X1 NAND2X1_910 ( .A(reg_hf__abc_3798_n115), .B(reg_hf__abc_3798_n114), .Y(reg_hf_value_11__FF_INPUT) );
	NOR2X1 NOR2X1_582 ( .A(reset), .B(reg_hf__abc_3798_n78), .Y(reg_hf__abc_3798_n117) );
	NAND2X1 NAND2X1_911 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n117), .Y(reg_hf__abc_3798_n118) );
	NAND2X1 NAND2X1_912 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n119) );
	NAND2X1 NAND2X1_913 ( .A(reg_hf__abc_3798_n119), .B(reg_hf__abc_3798_n118), .Y(reg_hf_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_583 ( .A(reset), .B(reg_hf__abc_3798_n80_1), .Y(reg_hf__abc_3798_n121) );
	NAND2X1 NAND2X1_914 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n121), .Y(reg_hf__abc_3798_n122) );
	NAND2X1 NAND2X1_915 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n123) );
	NAND2X1 NAND2X1_916 ( .A(reg_hf__abc_3798_n123), .B(reg_hf__abc_3798_n122), .Y(reg_hf__abc_3798_n50) );
	NOR2X1 NOR2X1_584 ( .A(reset), .B(reg_hf__abc_3798_n82_1), .Y(reg_hf__abc_3798_n125) );
	NAND2X1 NAND2X1_917 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n125), .Y(reg_hf__abc_3798_n126) );
	NAND2X1 NAND2X1_918 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n127) );
	NAND2X1 NAND2X1_919 ( .A(reg_hf__abc_3798_n127), .B(reg_hf__abc_3798_n126), .Y(reg_hf__abc_3798_n53) );
	NOR2X1 NOR2X1_585 ( .A(reset), .B(reg_hf__abc_3798_n84_1), .Y(reg_hf__abc_3798_n129) );
	NAND2X1 NAND2X1_920 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n129), .Y(reg_hf__abc_3798_n130) );
	NAND2X1 NAND2X1_921 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n131) );
	NAND2X1 NAND2X1_922 ( .A(reg_hf__abc_3798_n131), .B(reg_hf__abc_3798_n130), .Y(reg_hf__abc_3798_n56) );
	NOR2X1 NOR2X1_586 ( .A(reset), .B(reg_hf__abc_3798_n86), .Y(reg_hf__abc_3798_n133) );
	NAND2X1 NAND2X1_923 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n133), .Y(reg_hf__abc_3798_n134) );
	NAND2X1 NAND2X1_924 ( .A(reset), .B(vdd), .Y(reg_hf__abc_3798_n135) );
	NAND2X1 NAND2X1_925 ( .A(reg_hf__abc_3798_n135), .B(reg_hf__abc_3798_n134), .Y(reg_hf__abc_3798_n59) );
	NOR2X1 NOR2X1_587 ( .A(reset), .B(reg_hf__abc_3798_n88), .Y(reg_hf__abc_3798_n137) );
	NAND2X1 NAND2X1_926 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n137), .Y(reg_hf__abc_3798_n138) );
	NAND2X1 NAND2X1_927 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n139) );
	NAND2X1 NAND2X1_928 ( .A(reg_hf__abc_3798_n139), .B(reg_hf__abc_3798_n138), .Y(reg_hf__abc_3798_n62) );
	NOR2X1 NOR2X1_588 ( .A(reset), .B(reg_hf__abc_3798_n90), .Y(reg_hf__abc_3798_n141) );
	NAND2X1 NAND2X1_929 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n141), .Y(reg_hf__abc_3798_n142) );
	NAND2X1 NAND2X1_930 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n143) );
	NAND2X1 NAND2X1_931 ( .A(reg_hf__abc_3798_n143), .B(reg_hf__abc_3798_n142), .Y(reg_hf__abc_3798_n65) );
	NOR2X1 NOR2X1_589 ( .A(reset), .B(reg_hf__abc_3798_n92), .Y(reg_hf__abc_3798_n145) );
	NAND2X1 NAND2X1_932 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n145), .Y(reg_hf__abc_3798_n146) );
	NAND2X1 NAND2X1_933 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n147) );
	NAND2X1 NAND2X1_934 ( .A(reg_hf__abc_3798_n147), .B(reg_hf__abc_3798_n146), .Y(reg_hf__abc_3798_n68) );
	NOR2X1 NOR2X1_590 ( .A(reset), .B(reg_hf__abc_3798_n94), .Y(reg_hf__abc_3798_n149) );
	NAND2X1 NAND2X1_935 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n149), .Y(reg_hf__abc_3798_n150) );
	NAND2X1 NAND2X1_936 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n151) );
	NAND2X1 NAND2X1_937 ( .A(reg_hf__abc_3798_n151), .B(reg_hf__abc_3798_n150), .Y(reg_hf_value_2__FF_INPUT) );
	NOR2X1 NOR2X1_591 ( .A(reset), .B(reg_hf__abc_3798_n96), .Y(reg_hf__abc_3798_n153) );
	NAND2X1 NAND2X1_938 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n153), .Y(reg_hf__abc_3798_n154) );
	NAND2X1 NAND2X1_939 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n155) );
	NAND2X1 NAND2X1_940 ( .A(reg_hf__abc_3798_n155), .B(reg_hf__abc_3798_n154), .Y(reg_hf_value_1__FF_INPUT) );
	NOR2X1 NOR2X1_592 ( .A(reset), .B(reg_hf__abc_3798_n98), .Y(reg_hf__abc_3798_n157) );
	NAND2X1 NAND2X1_941 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n157), .Y(reg_hf__abc_3798_n158) );
	NAND2X1 NAND2X1_942 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n159) );
	NAND2X1 NAND2X1_943 ( .A(reg_hf__abc_3798_n159), .B(reg_hf__abc_3798_n158), .Y(reg_hf_value_0__FF_INPUT) );
	INVX1 INVX1_220 ( .A(reg_hf_value_15_), .Y(reg_hf__abc_3798_n161) );
	NOR2X1 NOR2X1_593 ( .A(reset), .B(reg_hf__abc_3798_n161), .Y(reg_hf__abc_3798_n162) );
	NAND2X1 NAND2X1_944 ( .A(reg_hf__abc_3798_n100), .B(reg_hf__abc_3798_n162), .Y(reg_hf__abc_3798_n163) );
	NAND2X1 NAND2X1_945 ( .A(reset), .B(gnd), .Y(reg_hf__abc_3798_n164) );
	NAND2X1 NAND2X1_946 ( .A(reg_hf__abc_3798_n164), .B(reg_hf__abc_3798_n163), .Y(reg_hf_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_594 ( .A(reg_hf__abc_3798_n161), .B(reg_hf__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_146 ( .CLK(clk), .D(reg_hf_value_0__FF_INPUT), .Q(reg_hf_value_0_) );
	DFFPOSX1 DFFPOSX1_147 ( .CLK(clk), .D(reg_hf_value_1__FF_INPUT), .Q(reg_hf_value_1_) );
	DFFPOSX1 DFFPOSX1_148 ( .CLK(clk), .D(reg_hf_value_2__FF_INPUT), .Q(reg_hf_value_2_) );
	DFFPOSX1 DFFPOSX1_149 ( .CLK(clk), .D(reg_hf__abc_3798_n68), .Q(reg_hf_value_3_) );
	DFFPOSX1 DFFPOSX1_150 ( .CLK(clk), .D(reg_hf__abc_3798_n65), .Q(reg_hf_value_4_) );
	DFFPOSX1 DFFPOSX1_151 ( .CLK(clk), .D(reg_hf__abc_3798_n62), .Q(reg_hf_value_5_) );
	DFFPOSX1 DFFPOSX1_152 ( .CLK(clk), .D(reg_hf__abc_3798_n59), .Q(reg_hf_value_6_) );
	DFFPOSX1 DFFPOSX1_153 ( .CLK(clk), .D(reg_hf__abc_3798_n56), .Q(reg_hf_value_7_) );
	DFFPOSX1 DFFPOSX1_154 ( .CLK(clk), .D(reg_hf__abc_3798_n53), .Q(reg_hf_value_8_) );
	DFFPOSX1 DFFPOSX1_155 ( .CLK(clk), .D(reg_hf__abc_3798_n50), .Q(reg_hf_value_9_) );
	DFFPOSX1 DFFPOSX1_156 ( .CLK(clk), .D(reg_hf_value_10__FF_INPUT), .Q(reg_hf_value_10_) );
	DFFPOSX1 DFFPOSX1_157 ( .CLK(clk), .D(reg_hf_value_11__FF_INPUT), .Q(reg_hf_value_11_) );
	DFFPOSX1 DFFPOSX1_158 ( .CLK(clk), .D(reg_hf_value_12__FF_INPUT), .Q(reg_hf_value_12_) );
	DFFPOSX1 DFFPOSX1_159 ( .CLK(clk), .D(reg_hf_value_13__FF_INPUT), .Q(reg_hf_value_13_) );
	DFFPOSX1 DFFPOSX1_160 ( .CLK(clk), .D(reg_hf_value_14__FF_INPUT), .Q(reg_hf_value_14_) );
	DFFPOSX1 DFFPOSX1_161 ( .CLK(clk), .D(reg_hf_value_15__FF_INPUT), .Q(reg_hf_value_15_) );
	INVX1 INVX1_221 ( .A(reg_hv_value_14_), .Y(reg_hv__abc_3798_n68_1) );
	INVX1 INVX1_222 ( .A(we), .Y(reg_hv__abc_3798_n69) );
	NAND2X1 NAND2X1_947 ( .A(addr_hv), .B(reg_hv__abc_3798_n69), .Y(reg_hv__abc_3798_n70_1) );
	NOR2X1 NOR2X1_595 ( .A(reg_hv__abc_3798_n68_1), .B(reg_hv__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_223 ( .A(reg_hv_value_13_), .Y(reg_hv__abc_3798_n72) );
	NOR2X1 NOR2X1_596 ( .A(reg_hv__abc_3798_n72), .B(reg_hv__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_224 ( .A(reg_hv_value_12_), .Y(reg_hv__abc_3798_n74_1) );
	NOR2X1 NOR2X1_597 ( .A(reg_hv__abc_3798_n74_1), .B(reg_hv__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_225 ( .A(reg_hv_value_11_), .Y(reg_hv__abc_3798_n76_1) );
	NOR2X1 NOR2X1_598 ( .A(reg_hv__abc_3798_n76_1), .B(reg_hv__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_226 ( .A(reg_hv_value_10_), .Y(reg_hv__abc_3798_n78) );
	NOR2X1 NOR2X1_599 ( .A(reg_hv__abc_3798_n78), .B(reg_hv__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_227 ( .A(reg_hv_value_9_), .Y(reg_hv__abc_3798_n80_1) );
	NOR2X1 NOR2X1_600 ( .A(reg_hv__abc_3798_n80_1), .B(reg_hv__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_228 ( .A(reg_hv_value_8_), .Y(reg_hv__abc_3798_n82_1) );
	NOR2X1 NOR2X1_601 ( .A(reg_hv__abc_3798_n82_1), .B(reg_hv__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_229 ( .A(reg_hv_value_7_), .Y(reg_hv__abc_3798_n84_1) );
	NOR2X1 NOR2X1_602 ( .A(reg_hv__abc_3798_n84_1), .B(reg_hv__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_230 ( .A(reg_hv_value_6_), .Y(reg_hv__abc_3798_n86) );
	NOR2X1 NOR2X1_603 ( .A(reg_hv__abc_3798_n86), .B(reg_hv__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_231 ( .A(reg_hv_value_5_), .Y(reg_hv__abc_3798_n88) );
	NOR2X1 NOR2X1_604 ( .A(reg_hv__abc_3798_n88), .B(reg_hv__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_232 ( .A(reg_hv_value_4_), .Y(reg_hv__abc_3798_n90) );
	NOR2X1 NOR2X1_605 ( .A(reg_hv__abc_3798_n90), .B(reg_hv__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_233 ( .A(reg_hv_value_3_), .Y(reg_hv__abc_3798_n92) );
	NOR2X1 NOR2X1_606 ( .A(reg_hv__abc_3798_n92), .B(reg_hv__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_234 ( .A(reg_hv_value_2_), .Y(reg_hv__abc_3798_n94) );
	NOR2X1 NOR2X1_607 ( .A(reg_hv__abc_3798_n94), .B(reg_hv__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_235 ( .A(reg_hv_value_1_), .Y(reg_hv__abc_3798_n96) );
	NOR2X1 NOR2X1_608 ( .A(reg_hv__abc_3798_n96), .B(reg_hv__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_236 ( .A(reg_hv_value_0_), .Y(reg_hv__abc_3798_n98) );
	NOR2X1 NOR2X1_609 ( .A(reg_hv__abc_3798_n98), .B(reg_hv__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_948 ( .A(we), .B(addr_hv), .Y(reg_hv__abc_3798_n100) );
	NOR2X1 NOR2X1_610 ( .A(reset), .B(reg_hv__abc_3798_n68_1), .Y(reg_hv__abc_3798_n101) );
	NAND2X1 NAND2X1_949 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n101), .Y(reg_hv__abc_3798_n102) );
	NAND2X1 NAND2X1_950 ( .A(gnd), .B(reset), .Y(reg_hv__abc_3798_n103) );
	NAND2X1 NAND2X1_951 ( .A(reg_hv__abc_3798_n103), .B(reg_hv__abc_3798_n102), .Y(reg_hv__abc_3798_n35) );
	NOR2X1 NOR2X1_611 ( .A(reset), .B(reg_hv__abc_3798_n72), .Y(reg_hv__abc_3798_n105) );
	NAND2X1 NAND2X1_952 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n105), .Y(reg_hv__abc_3798_n106) );
	NAND2X1 NAND2X1_953 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n107) );
	NAND2X1 NAND2X1_954 ( .A(reg_hv__abc_3798_n107), .B(reg_hv__abc_3798_n106), .Y(reg_hv__abc_3798_n38) );
	NOR2X1 NOR2X1_612 ( .A(reset), .B(reg_hv__abc_3798_n74_1), .Y(reg_hv__abc_3798_n109) );
	NAND2X1 NAND2X1_955 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n109), .Y(reg_hv__abc_3798_n110) );
	NAND2X1 NAND2X1_956 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n111) );
	NAND2X1 NAND2X1_957 ( .A(reg_hv__abc_3798_n111), .B(reg_hv__abc_3798_n110), .Y(reg_hv__abc_3798_n41) );
	NOR2X1 NOR2X1_613 ( .A(reset), .B(reg_hv__abc_3798_n76_1), .Y(reg_hv__abc_3798_n113) );
	NAND2X1 NAND2X1_958 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n113), .Y(reg_hv__abc_3798_n114) );
	NAND2X1 NAND2X1_959 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n115) );
	NAND2X1 NAND2X1_960 ( .A(reg_hv__abc_3798_n115), .B(reg_hv__abc_3798_n114), .Y(reg_hv__abc_3798_n44) );
	NOR2X1 NOR2X1_614 ( .A(reset), .B(reg_hv__abc_3798_n78), .Y(reg_hv__abc_3798_n117) );
	NAND2X1 NAND2X1_961 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n117), .Y(reg_hv__abc_3798_n118) );
	NAND2X1 NAND2X1_962 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n119) );
	NAND2X1 NAND2X1_963 ( .A(reg_hv__abc_3798_n119), .B(reg_hv__abc_3798_n118), .Y(reg_hv__abc_3798_n47) );
	NOR2X1 NOR2X1_615 ( .A(reset), .B(reg_hv__abc_3798_n80_1), .Y(reg_hv__abc_3798_n121) );
	NAND2X1 NAND2X1_964 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n121), .Y(reg_hv__abc_3798_n122) );
	NAND2X1 NAND2X1_965 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n123) );
	NAND2X1 NAND2X1_966 ( .A(reg_hv__abc_3798_n123), .B(reg_hv__abc_3798_n122), .Y(reg_hv__abc_3798_n50) );
	NOR2X1 NOR2X1_616 ( .A(reset), .B(reg_hv__abc_3798_n82_1), .Y(reg_hv__abc_3798_n125) );
	NAND2X1 NAND2X1_967 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n125), .Y(reg_hv__abc_3798_n126) );
	NAND2X1 NAND2X1_968 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n127) );
	NAND2X1 NAND2X1_969 ( .A(reg_hv__abc_3798_n127), .B(reg_hv__abc_3798_n126), .Y(reg_hv__abc_3798_n53) );
	NOR2X1 NOR2X1_617 ( .A(reset), .B(reg_hv__abc_3798_n84_1), .Y(reg_hv__abc_3798_n129) );
	NAND2X1 NAND2X1_970 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n129), .Y(reg_hv__abc_3798_n130) );
	NAND2X1 NAND2X1_971 ( .A(reset), .B(vdd), .Y(reg_hv__abc_3798_n131) );
	NAND2X1 NAND2X1_972 ( .A(reg_hv__abc_3798_n131), .B(reg_hv__abc_3798_n130), .Y(reg_hv__abc_3798_n56) );
	NOR2X1 NOR2X1_618 ( .A(reset), .B(reg_hv__abc_3798_n86), .Y(reg_hv__abc_3798_n133) );
	NAND2X1 NAND2X1_973 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n133), .Y(reg_hv__abc_3798_n134) );
	NAND2X1 NAND2X1_974 ( .A(reset), .B(vdd), .Y(reg_hv__abc_3798_n135) );
	NAND2X1 NAND2X1_975 ( .A(reg_hv__abc_3798_n135), .B(reg_hv__abc_3798_n134), .Y(reg_hv__abc_3798_n59) );
	NOR2X1 NOR2X1_619 ( .A(reset), .B(reg_hv__abc_3798_n88), .Y(reg_hv__abc_3798_n137) );
	NAND2X1 NAND2X1_976 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n137), .Y(reg_hv__abc_3798_n138) );
	NAND2X1 NAND2X1_977 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n139) );
	NAND2X1 NAND2X1_978 ( .A(reg_hv__abc_3798_n139), .B(reg_hv__abc_3798_n138), .Y(reg_hv__abc_3798_n62) );
	NOR2X1 NOR2X1_620 ( .A(reset), .B(reg_hv__abc_3798_n90), .Y(reg_hv__abc_3798_n141) );
	NAND2X1 NAND2X1_979 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n141), .Y(reg_hv__abc_3798_n142) );
	NAND2X1 NAND2X1_980 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n143) );
	NAND2X1 NAND2X1_981 ( .A(reg_hv__abc_3798_n143), .B(reg_hv__abc_3798_n142), .Y(reg_hv__abc_3798_n65) );
	NOR2X1 NOR2X1_621 ( .A(reset), .B(reg_hv__abc_3798_n92), .Y(reg_hv__abc_3798_n145) );
	NAND2X1 NAND2X1_982 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n145), .Y(reg_hv__abc_3798_n146) );
	NAND2X1 NAND2X1_983 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n147) );
	NAND2X1 NAND2X1_984 ( .A(reg_hv__abc_3798_n147), .B(reg_hv__abc_3798_n146), .Y(reg_hv__abc_3798_n68) );
	NOR2X1 NOR2X1_622 ( .A(reset), .B(reg_hv__abc_3798_n94), .Y(reg_hv__abc_3798_n149) );
	NAND2X1 NAND2X1_985 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n149), .Y(reg_hv__abc_3798_n150) );
	NAND2X1 NAND2X1_986 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n151) );
	NAND2X1 NAND2X1_987 ( .A(reg_hv__abc_3798_n151), .B(reg_hv__abc_3798_n150), .Y(reg_hv__abc_3798_n71) );
	NOR2X1 NOR2X1_623 ( .A(reset), .B(reg_hv__abc_3798_n96), .Y(reg_hv__abc_3798_n153) );
	NAND2X1 NAND2X1_988 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n153), .Y(reg_hv__abc_3798_n154) );
	NAND2X1 NAND2X1_989 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n155) );
	NAND2X1 NAND2X1_990 ( .A(reg_hv__abc_3798_n155), .B(reg_hv__abc_3798_n154), .Y(reg_hv__abc_3798_n74) );
	NOR2X1 NOR2X1_624 ( .A(reset), .B(reg_hv__abc_3798_n98), .Y(reg_hv__abc_3798_n157) );
	NAND2X1 NAND2X1_991 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n157), .Y(reg_hv__abc_3798_n158) );
	NAND2X1 NAND2X1_992 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n159) );
	NAND2X1 NAND2X1_993 ( .A(reg_hv__abc_3798_n159), .B(reg_hv__abc_3798_n158), .Y(reg_hv__abc_3798_n77) );
	INVX1 INVX1_237 ( .A(reg_hv_value_15_), .Y(reg_hv__abc_3798_n161) );
	NOR2X1 NOR2X1_625 ( .A(reset), .B(reg_hv__abc_3798_n161), .Y(reg_hv__abc_3798_n162) );
	NAND2X1 NAND2X1_994 ( .A(reg_hv__abc_3798_n100), .B(reg_hv__abc_3798_n162), .Y(reg_hv__abc_3798_n163) );
	NAND2X1 NAND2X1_995 ( .A(reset), .B(gnd), .Y(reg_hv__abc_3798_n164) );
	NAND2X1 NAND2X1_996 ( .A(reg_hv__abc_3798_n164), .B(reg_hv__abc_3798_n163), .Y(reg_hv__abc_3798_n81) );
	NOR2X1 NOR2X1_626 ( .A(reg_hv__abc_3798_n161), .B(reg_hv__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_162 ( .CLK(clk), .D(reg_hv__abc_3798_n77), .Q(reg_hv_value_0_) );
	DFFPOSX1 DFFPOSX1_163 ( .CLK(clk), .D(reg_hv__abc_3798_n74), .Q(reg_hv_value_1_) );
	DFFPOSX1 DFFPOSX1_164 ( .CLK(clk), .D(reg_hv__abc_3798_n71), .Q(reg_hv_value_2_) );
	DFFPOSX1 DFFPOSX1_165 ( .CLK(clk), .D(reg_hv__abc_3798_n68), .Q(reg_hv_value_3_) );
	DFFPOSX1 DFFPOSX1_166 ( .CLK(clk), .D(reg_hv__abc_3798_n65), .Q(reg_hv_value_4_) );
	DFFPOSX1 DFFPOSX1_167 ( .CLK(clk), .D(reg_hv__abc_3798_n62), .Q(reg_hv_value_5_) );
	DFFPOSX1 DFFPOSX1_168 ( .CLK(clk), .D(reg_hv__abc_3798_n59), .Q(reg_hv_value_6_) );
	DFFPOSX1 DFFPOSX1_169 ( .CLK(clk), .D(reg_hv__abc_3798_n56), .Q(reg_hv_value_7_) );
	DFFPOSX1 DFFPOSX1_170 ( .CLK(clk), .D(reg_hv__abc_3798_n53), .Q(reg_hv_value_8_) );
	DFFPOSX1 DFFPOSX1_171 ( .CLK(clk), .D(reg_hv__abc_3798_n50), .Q(reg_hv_value_9_) );
	DFFPOSX1 DFFPOSX1_172 ( .CLK(clk), .D(reg_hv__abc_3798_n47), .Q(reg_hv_value_10_) );
	DFFPOSX1 DFFPOSX1_173 ( .CLK(clk), .D(reg_hv__abc_3798_n44), .Q(reg_hv_value_11_) );
	DFFPOSX1 DFFPOSX1_174 ( .CLK(clk), .D(reg_hv__abc_3798_n41), .Q(reg_hv_value_12_) );
	DFFPOSX1 DFFPOSX1_175 ( .CLK(clk), .D(reg_hv__abc_3798_n38), .Q(reg_hv_value_13_) );
	DFFPOSX1 DFFPOSX1_176 ( .CLK(clk), .D(reg_hv__abc_3798_n35), .Q(reg_hv_value_14_) );
	DFFPOSX1 DFFPOSX1_177 ( .CLK(clk), .D(reg_hv__abc_3798_n81), .Q(reg_hv_value_15_) );
	INVX1 INVX1_238 ( .A(reg_ic_value_14_), .Y(reg_ic__abc_3798_n68_1) );
	INVX1 INVX1_239 ( .A(we), .Y(reg_ic__abc_3798_n69) );
	NAND2X1 NAND2X1_997 ( .A(addr_ic), .B(reg_ic__abc_3798_n69), .Y(reg_ic__abc_3798_n70_1) );
	NOR2X1 NOR2X1_627 ( .A(reg_ic__abc_3798_n68_1), .B(reg_ic__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_240 ( .A(reg_ic_value_13_), .Y(reg_ic__abc_3798_n72) );
	NOR2X1 NOR2X1_628 ( .A(reg_ic__abc_3798_n72), .B(reg_ic__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_241 ( .A(reg_ic_value_12_), .Y(reg_ic__abc_3798_n74_1) );
	NOR2X1 NOR2X1_629 ( .A(reg_ic__abc_3798_n74_1), .B(reg_ic__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_242 ( .A(reg_ic_value_11_), .Y(reg_ic__abc_3798_n76_1) );
	NOR2X1 NOR2X1_630 ( .A(reg_ic__abc_3798_n76_1), .B(reg_ic__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_243 ( .A(reg_ic_value_10_), .Y(reg_ic__abc_3798_n78) );
	NOR2X1 NOR2X1_631 ( .A(reg_ic__abc_3798_n78), .B(reg_ic__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_244 ( .A(reg_ic_value_9_), .Y(reg_ic__abc_3798_n80_1) );
	NOR2X1 NOR2X1_632 ( .A(reg_ic__abc_3798_n80_1), .B(reg_ic__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_245 ( .A(reg_ic_value_8_), .Y(reg_ic__abc_3798_n82_1) );
	NOR2X1 NOR2X1_633 ( .A(reg_ic__abc_3798_n82_1), .B(reg_ic__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_246 ( .A(reg_ic_value_7_), .Y(reg_ic__abc_3798_n84_1) );
	NOR2X1 NOR2X1_634 ( .A(reg_ic__abc_3798_n84_1), .B(reg_ic__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_247 ( .A(reg_ic_value_6_), .Y(reg_ic__abc_3798_n86) );
	NOR2X1 NOR2X1_635 ( .A(reg_ic__abc_3798_n86), .B(reg_ic__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_248 ( .A(reg_ic_value_5_), .Y(reg_ic__abc_3798_n88) );
	NOR2X1 NOR2X1_636 ( .A(reg_ic__abc_3798_n88), .B(reg_ic__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_249 ( .A(reg_ic_value_4_), .Y(reg_ic__abc_3798_n90) );
	NOR2X1 NOR2X1_637 ( .A(reg_ic__abc_3798_n90), .B(reg_ic__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_250 ( .A(reg_ic_value_3_), .Y(reg_ic__abc_3798_n92) );
	NOR2X1 NOR2X1_638 ( .A(reg_ic__abc_3798_n92), .B(reg_ic__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_251 ( .A(reg_ic_value_2_), .Y(reg_ic__abc_3798_n94) );
	NOR2X1 NOR2X1_639 ( .A(reg_ic__abc_3798_n94), .B(reg_ic__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_252 ( .A(reg_ic_value_1_), .Y(reg_ic__abc_3798_n96) );
	NOR2X1 NOR2X1_640 ( .A(reg_ic__abc_3798_n96), .B(reg_ic__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_253 ( .A(reg_ic_value_0_), .Y(reg_ic__abc_3798_n98) );
	NOR2X1 NOR2X1_641 ( .A(reg_ic__abc_3798_n98), .B(reg_ic__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_998 ( .A(we), .B(addr_ic), .Y(reg_ic__abc_3798_n100) );
	NOR2X1 NOR2X1_642 ( .A(reset), .B(reg_ic__abc_3798_n68_1), .Y(reg_ic__abc_3798_n101) );
	NAND2X1 NAND2X1_999 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n101), .Y(reg_ic__abc_3798_n102) );
	NAND2X1 NAND2X1_1000 ( .A(gnd), .B(reset), .Y(reg_ic__abc_3798_n103) );
	NAND2X1 NAND2X1_1001 ( .A(reg_ic__abc_3798_n103), .B(reg_ic__abc_3798_n102), .Y(reg_ic__abc_3798_n35) );
	NOR2X1 NOR2X1_643 ( .A(reset), .B(reg_ic__abc_3798_n72), .Y(reg_ic__abc_3798_n105) );
	NAND2X1 NAND2X1_1002 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n105), .Y(reg_ic__abc_3798_n106) );
	NAND2X1 NAND2X1_1003 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n107) );
	NAND2X1 NAND2X1_1004 ( .A(reg_ic__abc_3798_n107), .B(reg_ic__abc_3798_n106), .Y(reg_ic__abc_3798_n38) );
	NOR2X1 NOR2X1_644 ( .A(reset), .B(reg_ic__abc_3798_n74_1), .Y(reg_ic__abc_3798_n109) );
	NAND2X1 NAND2X1_1005 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n109), .Y(reg_ic__abc_3798_n110) );
	NAND2X1 NAND2X1_1006 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n111) );
	NAND2X1 NAND2X1_1007 ( .A(reg_ic__abc_3798_n111), .B(reg_ic__abc_3798_n110), .Y(reg_ic__abc_3798_n41) );
	NOR2X1 NOR2X1_645 ( .A(reset), .B(reg_ic__abc_3798_n76_1), .Y(reg_ic__abc_3798_n113) );
	NAND2X1 NAND2X1_1008 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n113), .Y(reg_ic__abc_3798_n114) );
	NAND2X1 NAND2X1_1009 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n115) );
	NAND2X1 NAND2X1_1010 ( .A(reg_ic__abc_3798_n115), .B(reg_ic__abc_3798_n114), .Y(reg_ic__abc_3798_n44) );
	NOR2X1 NOR2X1_646 ( .A(reset), .B(reg_ic__abc_3798_n78), .Y(reg_ic__abc_3798_n117) );
	NAND2X1 NAND2X1_1011 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n117), .Y(reg_ic__abc_3798_n118) );
	NAND2X1 NAND2X1_1012 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n119) );
	NAND2X1 NAND2X1_1013 ( .A(reg_ic__abc_3798_n119), .B(reg_ic__abc_3798_n118), .Y(reg_ic__abc_3798_n47) );
	NOR2X1 NOR2X1_647 ( .A(reset), .B(reg_ic__abc_3798_n80_1), .Y(reg_ic__abc_3798_n121) );
	NAND2X1 NAND2X1_1014 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n121), .Y(reg_ic__abc_3798_n122) );
	NAND2X1 NAND2X1_1015 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n123) );
	NAND2X1 NAND2X1_1016 ( .A(reg_ic__abc_3798_n123), .B(reg_ic__abc_3798_n122), .Y(reg_ic__abc_3798_n50) );
	NOR2X1 NOR2X1_648 ( .A(reset), .B(reg_ic__abc_3798_n82_1), .Y(reg_ic__abc_3798_n125) );
	NAND2X1 NAND2X1_1017 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n125), .Y(reg_ic__abc_3798_n126) );
	NAND2X1 NAND2X1_1018 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n127) );
	NAND2X1 NAND2X1_1019 ( .A(reg_ic__abc_3798_n127), .B(reg_ic__abc_3798_n126), .Y(reg_ic__abc_3798_n53) );
	NOR2X1 NOR2X1_649 ( .A(reset), .B(reg_ic__abc_3798_n84_1), .Y(reg_ic__abc_3798_n129) );
	NAND2X1 NAND2X1_1020 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n129), .Y(reg_ic__abc_3798_n130) );
	NAND2X1 NAND2X1_1021 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n131) );
	NAND2X1 NAND2X1_1022 ( .A(reg_ic__abc_3798_n131), .B(reg_ic__abc_3798_n130), .Y(reg_ic__abc_3798_n56) );
	NOR2X1 NOR2X1_650 ( .A(reset), .B(reg_ic__abc_3798_n86), .Y(reg_ic__abc_3798_n133) );
	NAND2X1 NAND2X1_1023 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n133), .Y(reg_ic__abc_3798_n134) );
	NAND2X1 NAND2X1_1024 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n135) );
	NAND2X1 NAND2X1_1025 ( .A(reg_ic__abc_3798_n135), .B(reg_ic__abc_3798_n134), .Y(reg_ic__abc_3798_n59) );
	NOR2X1 NOR2X1_651 ( .A(reset), .B(reg_ic__abc_3798_n88), .Y(reg_ic__abc_3798_n137) );
	NAND2X1 NAND2X1_1026 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n137), .Y(reg_ic__abc_3798_n138) );
	NAND2X1 NAND2X1_1027 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n139) );
	NAND2X1 NAND2X1_1028 ( .A(reg_ic__abc_3798_n139), .B(reg_ic__abc_3798_n138), .Y(reg_ic__abc_3798_n62) );
	NOR2X1 NOR2X1_652 ( .A(reset), .B(reg_ic__abc_3798_n90), .Y(reg_ic__abc_3798_n141) );
	NAND2X1 NAND2X1_1029 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n141), .Y(reg_ic__abc_3798_n142) );
	NAND2X1 NAND2X1_1030 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n143) );
	NAND2X1 NAND2X1_1031 ( .A(reg_ic__abc_3798_n143), .B(reg_ic__abc_3798_n142), .Y(reg_ic__abc_3798_n65) );
	NOR2X1 NOR2X1_653 ( .A(reset), .B(reg_ic__abc_3798_n92), .Y(reg_ic__abc_3798_n145) );
	NAND2X1 NAND2X1_1032 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n145), .Y(reg_ic__abc_3798_n146) );
	NAND2X1 NAND2X1_1033 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n147) );
	NAND2X1 NAND2X1_1034 ( .A(reg_ic__abc_3798_n147), .B(reg_ic__abc_3798_n146), .Y(reg_ic__abc_3798_n68) );
	NOR2X1 NOR2X1_654 ( .A(reset), .B(reg_ic__abc_3798_n94), .Y(reg_ic__abc_3798_n149) );
	NAND2X1 NAND2X1_1035 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n149), .Y(reg_ic__abc_3798_n150) );
	NAND2X1 NAND2X1_1036 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n151) );
	NAND2X1 NAND2X1_1037 ( .A(reg_ic__abc_3798_n151), .B(reg_ic__abc_3798_n150), .Y(reg_ic__abc_3798_n71) );
	NOR2X1 NOR2X1_655 ( .A(reset), .B(reg_ic__abc_3798_n96), .Y(reg_ic__abc_3798_n153) );
	NAND2X1 NAND2X1_1038 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n153), .Y(reg_ic__abc_3798_n154) );
	NAND2X1 NAND2X1_1039 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n155) );
	NAND2X1 NAND2X1_1040 ( .A(reg_ic__abc_3798_n155), .B(reg_ic__abc_3798_n154), .Y(reg_ic__abc_3798_n74) );
	NOR2X1 NOR2X1_656 ( .A(reset), .B(reg_ic__abc_3798_n98), .Y(reg_ic__abc_3798_n157) );
	NAND2X1 NAND2X1_1041 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n157), .Y(reg_ic__abc_3798_n158) );
	NAND2X1 NAND2X1_1042 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n159) );
	NAND2X1 NAND2X1_1043 ( .A(reg_ic__abc_3798_n159), .B(reg_ic__abc_3798_n158), .Y(reg_ic__abc_3798_n77) );
	INVX1 INVX1_254 ( .A(reg_ic_value_15_), .Y(reg_ic__abc_3798_n161) );
	NOR2X1 NOR2X1_657 ( .A(reset), .B(reg_ic__abc_3798_n161), .Y(reg_ic__abc_3798_n162) );
	NAND2X1 NAND2X1_1044 ( .A(reg_ic__abc_3798_n100), .B(reg_ic__abc_3798_n162), .Y(reg_ic__abc_3798_n163) );
	NAND2X1 NAND2X1_1045 ( .A(reset), .B(gnd), .Y(reg_ic__abc_3798_n164) );
	NAND2X1 NAND2X1_1046 ( .A(reg_ic__abc_3798_n164), .B(reg_ic__abc_3798_n163), .Y(reg_ic__abc_3798_n81) );
	NOR2X1 NOR2X1_658 ( .A(reg_ic__abc_3798_n161), .B(reg_ic__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_178 ( .CLK(clk), .D(reg_ic__abc_3798_n77), .Q(reg_ic_value_0_) );
	DFFPOSX1 DFFPOSX1_179 ( .CLK(clk), .D(reg_ic__abc_3798_n74), .Q(reg_ic_value_1_) );
	DFFPOSX1 DFFPOSX1_180 ( .CLK(clk), .D(reg_ic__abc_3798_n71), .Q(reg_ic_value_2_) );
	DFFPOSX1 DFFPOSX1_181 ( .CLK(clk), .D(reg_ic__abc_3798_n68), .Q(reg_ic_value_3_) );
	DFFPOSX1 DFFPOSX1_182 ( .CLK(clk), .D(reg_ic__abc_3798_n65), .Q(reg_ic_value_4_) );
	DFFPOSX1 DFFPOSX1_183 ( .CLK(clk), .D(reg_ic__abc_3798_n62), .Q(reg_ic_value_5_) );
	DFFPOSX1 DFFPOSX1_184 ( .CLK(clk), .D(reg_ic__abc_3798_n59), .Q(reg_ic_value_6_) );
	DFFPOSX1 DFFPOSX1_185 ( .CLK(clk), .D(reg_ic__abc_3798_n56), .Q(reg_ic_value_7_) );
	DFFPOSX1 DFFPOSX1_186 ( .CLK(clk), .D(reg_ic__abc_3798_n53), .Q(reg_ic_value_8_) );
	DFFPOSX1 DFFPOSX1_187 ( .CLK(clk), .D(reg_ic__abc_3798_n50), .Q(reg_ic_value_9_) );
	DFFPOSX1 DFFPOSX1_188 ( .CLK(clk), .D(reg_ic__abc_3798_n47), .Q(reg_ic_value_10_) );
	DFFPOSX1 DFFPOSX1_189 ( .CLK(clk), .D(reg_ic__abc_3798_n44), .Q(reg_ic_value_11_) );
	DFFPOSX1 DFFPOSX1_190 ( .CLK(clk), .D(reg_ic__abc_3798_n41), .Q(reg_ic_value_12_) );
	DFFPOSX1 DFFPOSX1_191 ( .CLK(clk), .D(reg_ic__abc_3798_n38), .Q(reg_ic_value_13_) );
	DFFPOSX1 DFFPOSX1_192 ( .CLK(clk), .D(reg_ic__abc_3798_n35), .Q(reg_ic_value_14_) );
	DFFPOSX1 DFFPOSX1_193 ( .CLK(clk), .D(reg_ic__abc_3798_n81), .Q(reg_ic_value_15_) );
	INVX1 INVX1_255 ( .A(reg_ir_value_14_), .Y(reg_ir__abc_3798_n68_1) );
	INVX1 INVX1_256 ( .A(we), .Y(reg_ir__abc_3798_n69) );
	NAND2X1 NAND2X1_1047 ( .A(addr_ir), .B(reg_ir__abc_3798_n69), .Y(reg_ir__abc_3798_n70_1) );
	NOR2X1 NOR2X1_659 ( .A(reg_ir__abc_3798_n68_1), .B(reg_ir__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_257 ( .A(reg_ir_value_13_), .Y(reg_ir__abc_3798_n72) );
	NOR2X1 NOR2X1_660 ( .A(reg_ir__abc_3798_n72), .B(reg_ir__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_258 ( .A(reg_ir_value_12_), .Y(reg_ir__abc_3798_n74_1) );
	NOR2X1 NOR2X1_661 ( .A(reg_ir__abc_3798_n74_1), .B(reg_ir__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_259 ( .A(reg_ir_value_11_), .Y(reg_ir__abc_3798_n76_1) );
	NOR2X1 NOR2X1_662 ( .A(reg_ir__abc_3798_n76_1), .B(reg_ir__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_260 ( .A(reg_ir_value_10_), .Y(reg_ir__abc_3798_n78) );
	NOR2X1 NOR2X1_663 ( .A(reg_ir__abc_3798_n78), .B(reg_ir__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_261 ( .A(reg_ir_value_9_), .Y(reg_ir__abc_3798_n80_1) );
	NOR2X1 NOR2X1_664 ( .A(reg_ir__abc_3798_n80_1), .B(reg_ir__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_262 ( .A(reg_ir_value_8_), .Y(reg_ir__abc_3798_n82_1) );
	NOR2X1 NOR2X1_665 ( .A(reg_ir__abc_3798_n82_1), .B(reg_ir__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_263 ( .A(reg_ir_value_7_), .Y(reg_ir__abc_3798_n84_1) );
	NOR2X1 NOR2X1_666 ( .A(reg_ir__abc_3798_n84_1), .B(reg_ir__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_264 ( .A(reg_ir_value_6_), .Y(reg_ir__abc_3798_n86) );
	NOR2X1 NOR2X1_667 ( .A(reg_ir__abc_3798_n86), .B(reg_ir__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_265 ( .A(reg_ir_value_5_), .Y(reg_ir__abc_3798_n88) );
	NOR2X1 NOR2X1_668 ( .A(reg_ir__abc_3798_n88), .B(reg_ir__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_266 ( .A(reg_ir_value_4_), .Y(reg_ir__abc_3798_n90) );
	NOR2X1 NOR2X1_669 ( .A(reg_ir__abc_3798_n90), .B(reg_ir__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_267 ( .A(reg_ir_value_3_), .Y(reg_ir__abc_3798_n92) );
	NOR2X1 NOR2X1_670 ( .A(reg_ir__abc_3798_n92), .B(reg_ir__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_268 ( .A(reg_ir_value_2_), .Y(reg_ir__abc_3798_n94) );
	NOR2X1 NOR2X1_671 ( .A(reg_ir__abc_3798_n94), .B(reg_ir__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_269 ( .A(reg_ir_value_1_), .Y(reg_ir__abc_3798_n96) );
	NOR2X1 NOR2X1_672 ( .A(reg_ir__abc_3798_n96), .B(reg_ir__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_270 ( .A(reg_ir_value_0_), .Y(reg_ir__abc_3798_n98) );
	NOR2X1 NOR2X1_673 ( .A(reg_ir__abc_3798_n98), .B(reg_ir__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1048 ( .A(we), .B(addr_ir), .Y(reg_ir__abc_3798_n100) );
	NOR2X1 NOR2X1_674 ( .A(reset), .B(reg_ir__abc_3798_n68_1), .Y(reg_ir__abc_3798_n101) );
	NAND2X1 NAND2X1_1049 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n101), .Y(reg_ir__abc_3798_n102) );
	NAND2X1 NAND2X1_1050 ( .A(gnd), .B(reset), .Y(reg_ir__abc_3798_n103) );
	NAND2X1 NAND2X1_1051 ( .A(reg_ir__abc_3798_n103), .B(reg_ir__abc_3798_n102), .Y(reg_ir_value_14__FF_INPUT) );
	NOR2X1 NOR2X1_675 ( .A(reset), .B(reg_ir__abc_3798_n72), .Y(reg_ir__abc_3798_n105) );
	NAND2X1 NAND2X1_1052 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n105), .Y(reg_ir__abc_3798_n106) );
	NAND2X1 NAND2X1_1053 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n107) );
	NAND2X1 NAND2X1_1054 ( .A(reg_ir__abc_3798_n107), .B(reg_ir__abc_3798_n106), .Y(reg_ir_value_13__FF_INPUT) );
	NOR2X1 NOR2X1_676 ( .A(reset), .B(reg_ir__abc_3798_n74_1), .Y(reg_ir__abc_3798_n109) );
	NAND2X1 NAND2X1_1055 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n109), .Y(reg_ir__abc_3798_n110) );
	NAND2X1 NAND2X1_1056 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n111) );
	NAND2X1 NAND2X1_1057 ( .A(reg_ir__abc_3798_n111), .B(reg_ir__abc_3798_n110), .Y(reg_ir_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_677 ( .A(reset), .B(reg_ir__abc_3798_n76_1), .Y(reg_ir__abc_3798_n113) );
	NAND2X1 NAND2X1_1058 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n113), .Y(reg_ir__abc_3798_n114) );
	NAND2X1 NAND2X1_1059 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n115) );
	NAND2X1 NAND2X1_1060 ( .A(reg_ir__abc_3798_n115), .B(reg_ir__abc_3798_n114), .Y(reg_ir_value_11__FF_INPUT) );
	NOR2X1 NOR2X1_678 ( .A(reset), .B(reg_ir__abc_3798_n78), .Y(reg_ir__abc_3798_n117) );
	NAND2X1 NAND2X1_1061 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n117), .Y(reg_ir__abc_3798_n118) );
	NAND2X1 NAND2X1_1062 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n119) );
	NAND2X1 NAND2X1_1063 ( .A(reg_ir__abc_3798_n119), .B(reg_ir__abc_3798_n118), .Y(reg_ir_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_679 ( .A(reset), .B(reg_ir__abc_3798_n80_1), .Y(reg_ir__abc_3798_n121) );
	NAND2X1 NAND2X1_1064 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n121), .Y(reg_ir__abc_3798_n122) );
	NAND2X1 NAND2X1_1065 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n123) );
	NAND2X1 NAND2X1_1066 ( .A(reg_ir__abc_3798_n123), .B(reg_ir__abc_3798_n122), .Y(reg_ir_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_680 ( .A(reset), .B(reg_ir__abc_3798_n82_1), .Y(reg_ir__abc_3798_n125) );
	NAND2X1 NAND2X1_1067 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n125), .Y(reg_ir__abc_3798_n126) );
	NAND2X1 NAND2X1_1068 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n127) );
	NAND2X1 NAND2X1_1069 ( .A(reg_ir__abc_3798_n127), .B(reg_ir__abc_3798_n126), .Y(reg_ir_value_8__FF_INPUT) );
	NOR2X1 NOR2X1_681 ( .A(reset), .B(reg_ir__abc_3798_n84_1), .Y(reg_ir__abc_3798_n129) );
	NAND2X1 NAND2X1_1070 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n129), .Y(reg_ir__abc_3798_n130) );
	NAND2X1 NAND2X1_1071 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n131) );
	NAND2X1 NAND2X1_1072 ( .A(reg_ir__abc_3798_n131), .B(reg_ir__abc_3798_n130), .Y(reg_ir_value_7__FF_INPUT) );
	NOR2X1 NOR2X1_682 ( .A(reset), .B(reg_ir__abc_3798_n86), .Y(reg_ir__abc_3798_n133) );
	NAND2X1 NAND2X1_1073 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n133), .Y(reg_ir__abc_3798_n134) );
	NAND2X1 NAND2X1_1074 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n135) );
	NAND2X1 NAND2X1_1075 ( .A(reg_ir__abc_3798_n135), .B(reg_ir__abc_3798_n134), .Y(reg_ir_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_683 ( .A(reset), .B(reg_ir__abc_3798_n88), .Y(reg_ir__abc_3798_n137) );
	NAND2X1 NAND2X1_1076 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n137), .Y(reg_ir__abc_3798_n138) );
	NAND2X1 NAND2X1_1077 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n139) );
	NAND2X1 NAND2X1_1078 ( .A(reg_ir__abc_3798_n139), .B(reg_ir__abc_3798_n138), .Y(reg_ir_value_5__FF_INPUT) );
	NOR2X1 NOR2X1_684 ( .A(reset), .B(reg_ir__abc_3798_n90), .Y(reg_ir__abc_3798_n141) );
	NAND2X1 NAND2X1_1079 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n141), .Y(reg_ir__abc_3798_n142) );
	NAND2X1 NAND2X1_1080 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n143) );
	NAND2X1 NAND2X1_1081 ( .A(reg_ir__abc_3798_n143), .B(reg_ir__abc_3798_n142), .Y(reg_ir_value_4__FF_INPUT) );
	NOR2X1 NOR2X1_685 ( .A(reset), .B(reg_ir__abc_3798_n92), .Y(reg_ir__abc_3798_n145) );
	NAND2X1 NAND2X1_1082 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n145), .Y(reg_ir__abc_3798_n146) );
	NAND2X1 NAND2X1_1083 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n147) );
	NAND2X1 NAND2X1_1084 ( .A(reg_ir__abc_3798_n147), .B(reg_ir__abc_3798_n146), .Y(reg_ir_value_3__FF_INPUT) );
	NOR2X1 NOR2X1_686 ( .A(reset), .B(reg_ir__abc_3798_n94), .Y(reg_ir__abc_3798_n149) );
	NAND2X1 NAND2X1_1085 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n149), .Y(reg_ir__abc_3798_n150) );
	NAND2X1 NAND2X1_1086 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n151) );
	NAND2X1 NAND2X1_1087 ( .A(reg_ir__abc_3798_n151), .B(reg_ir__abc_3798_n150), .Y(reg_ir_value_2__FF_INPUT) );
	NOR2X1 NOR2X1_687 ( .A(reset), .B(reg_ir__abc_3798_n96), .Y(reg_ir__abc_3798_n153) );
	NAND2X1 NAND2X1_1088 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n153), .Y(reg_ir__abc_3798_n154) );
	NAND2X1 NAND2X1_1089 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n155) );
	NAND2X1 NAND2X1_1090 ( .A(reg_ir__abc_3798_n155), .B(reg_ir__abc_3798_n154), .Y(reg_ir_value_1__FF_INPUT) );
	NOR2X1 NOR2X1_688 ( .A(reset), .B(reg_ir__abc_3798_n98), .Y(reg_ir__abc_3798_n157) );
	NAND2X1 NAND2X1_1091 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n157), .Y(reg_ir__abc_3798_n158) );
	NAND2X1 NAND2X1_1092 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n159) );
	NAND2X1 NAND2X1_1093 ( .A(reg_ir__abc_3798_n159), .B(reg_ir__abc_3798_n158), .Y(reg_ir_value_0__FF_INPUT) );
	INVX1 INVX1_271 ( .A(reg_ir_value_15_), .Y(reg_ir__abc_3798_n161) );
	NOR2X1 NOR2X1_689 ( .A(reset), .B(reg_ir__abc_3798_n161), .Y(reg_ir__abc_3798_n162) );
	NAND2X1 NAND2X1_1094 ( .A(reg_ir__abc_3798_n100), .B(reg_ir__abc_3798_n162), .Y(reg_ir__abc_3798_n163) );
	NAND2X1 NAND2X1_1095 ( .A(reset), .B(gnd), .Y(reg_ir__abc_3798_n164) );
	NAND2X1 NAND2X1_1096 ( .A(reg_ir__abc_3798_n164), .B(reg_ir__abc_3798_n163), .Y(reg_ir_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_690 ( .A(reg_ir__abc_3798_n161), .B(reg_ir__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_194 ( .CLK(clk), .D(reg_ir_value_0__FF_INPUT), .Q(reg_ir_value_0_) );
	DFFPOSX1 DFFPOSX1_195 ( .CLK(clk), .D(reg_ir_value_1__FF_INPUT), .Q(reg_ir_value_1_) );
	DFFPOSX1 DFFPOSX1_196 ( .CLK(clk), .D(reg_ir_value_2__FF_INPUT), .Q(reg_ir_value_2_) );
	DFFPOSX1 DFFPOSX1_197 ( .CLK(clk), .D(reg_ir_value_3__FF_INPUT), .Q(reg_ir_value_3_) );
	DFFPOSX1 DFFPOSX1_198 ( .CLK(clk), .D(reg_ir_value_4__FF_INPUT), .Q(reg_ir_value_4_) );
	DFFPOSX1 DFFPOSX1_199 ( .CLK(clk), .D(reg_ir_value_5__FF_INPUT), .Q(reg_ir_value_5_) );
	DFFPOSX1 DFFPOSX1_200 ( .CLK(clk), .D(reg_ir_value_6__FF_INPUT), .Q(reg_ir_value_6_) );
	DFFPOSX1 DFFPOSX1_201 ( .CLK(clk), .D(reg_ir_value_7__FF_INPUT), .Q(reg_ir_value_7_) );
	DFFPOSX1 DFFPOSX1_202 ( .CLK(clk), .D(reg_ir_value_8__FF_INPUT), .Q(reg_ir_value_8_) );
	DFFPOSX1 DFFPOSX1_203 ( .CLK(clk), .D(reg_ir_value_9__FF_INPUT), .Q(reg_ir_value_9_) );
	DFFPOSX1 DFFPOSX1_204 ( .CLK(clk), .D(reg_ir_value_10__FF_INPUT), .Q(reg_ir_value_10_) );
	DFFPOSX1 DFFPOSX1_205 ( .CLK(clk), .D(reg_ir_value_11__FF_INPUT), .Q(reg_ir_value_11_) );
	DFFPOSX1 DFFPOSX1_206 ( .CLK(clk), .D(reg_ir_value_12__FF_INPUT), .Q(reg_ir_value_12_) );
	DFFPOSX1 DFFPOSX1_207 ( .CLK(clk), .D(reg_ir_value_13__FF_INPUT), .Q(reg_ir_value_13_) );
	DFFPOSX1 DFFPOSX1_208 ( .CLK(clk), .D(reg_ir_value_14__FF_INPUT), .Q(reg_ir_value_14_) );
	DFFPOSX1 DFFPOSX1_209 ( .CLK(clk), .D(reg_ir_value_15__FF_INPUT), .Q(reg_ir_value_15_) );
	INVX1 INVX1_272 ( .A(reg_sh_value_14_), .Y(reg_sh__abc_3798_n68_1) );
	INVX1 INVX1_273 ( .A(we), .Y(reg_sh__abc_3798_n69) );
	NAND2X1 NAND2X1_1097 ( .A(addr_sh), .B(reg_sh__abc_3798_n69), .Y(reg_sh__abc_3798_n70_1) );
	NOR2X1 NOR2X1_691 ( .A(reg_sh__abc_3798_n68_1), .B(reg_sh__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_274 ( .A(reg_sh_value_13_), .Y(reg_sh__abc_3798_n72) );
	NOR2X1 NOR2X1_692 ( .A(reg_sh__abc_3798_n72), .B(reg_sh__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_275 ( .A(reg_sh_value_12_), .Y(reg_sh__abc_3798_n74_1) );
	NOR2X1 NOR2X1_693 ( .A(reg_sh__abc_3798_n74_1), .B(reg_sh__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_276 ( .A(reg_sh_value_11_), .Y(reg_sh__abc_3798_n76_1) );
	NOR2X1 NOR2X1_694 ( .A(reg_sh__abc_3798_n76_1), .B(reg_sh__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_277 ( .A(reg_sh_value_10_), .Y(reg_sh__abc_3798_n78) );
	NOR2X1 NOR2X1_695 ( .A(reg_sh__abc_3798_n78), .B(reg_sh__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_278 ( .A(reg_sh_value_9_), .Y(reg_sh__abc_3798_n80_1) );
	NOR2X1 NOR2X1_696 ( .A(reg_sh__abc_3798_n80_1), .B(reg_sh__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_279 ( .A(reg_sh_value_8_), .Y(reg_sh__abc_3798_n82_1) );
	NOR2X1 NOR2X1_697 ( .A(reg_sh__abc_3798_n82_1), .B(reg_sh__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_280 ( .A(reg_sh_value_7_), .Y(reg_sh__abc_3798_n84_1) );
	NOR2X1 NOR2X1_698 ( .A(reg_sh__abc_3798_n84_1), .B(reg_sh__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_281 ( .A(reg_sh_value_6_), .Y(reg_sh__abc_3798_n86) );
	NOR2X1 NOR2X1_699 ( .A(reg_sh__abc_3798_n86), .B(reg_sh__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_282 ( .A(reg_sh_value_5_), .Y(reg_sh__abc_3798_n88) );
	NOR2X1 NOR2X1_700 ( .A(reg_sh__abc_3798_n88), .B(reg_sh__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_283 ( .A(reg_sh_value_4_), .Y(reg_sh__abc_3798_n90) );
	NOR2X1 NOR2X1_701 ( .A(reg_sh__abc_3798_n90), .B(reg_sh__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_284 ( .A(reg_sh_value_3_), .Y(reg_sh__abc_3798_n92) );
	NOR2X1 NOR2X1_702 ( .A(reg_sh__abc_3798_n92), .B(reg_sh__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_285 ( .A(reg_sh_value_2_), .Y(reg_sh__abc_3798_n94) );
	NOR2X1 NOR2X1_703 ( .A(reg_sh__abc_3798_n94), .B(reg_sh__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_286 ( .A(reg_sh_value_1_), .Y(reg_sh__abc_3798_n96) );
	NOR2X1 NOR2X1_704 ( .A(reg_sh__abc_3798_n96), .B(reg_sh__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_287 ( .A(reg_sh_value_0_), .Y(reg_sh__abc_3798_n98) );
	NOR2X1 NOR2X1_705 ( .A(reg_sh__abc_3798_n98), .B(reg_sh__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1098 ( .A(we), .B(addr_sh), .Y(reg_sh__abc_3798_n100) );
	NOR2X1 NOR2X1_706 ( .A(reset), .B(reg_sh__abc_3798_n68_1), .Y(reg_sh__abc_3798_n101) );
	NAND2X1 NAND2X1_1099 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n101), .Y(reg_sh__abc_3798_n102) );
	NAND2X1 NAND2X1_1100 ( .A(gnd), .B(reset), .Y(reg_sh__abc_3798_n103) );
	NAND2X1 NAND2X1_1101 ( .A(reg_sh__abc_3798_n103), .B(reg_sh__abc_3798_n102), .Y(reg_sh_value_14__FF_INPUT) );
	NOR2X1 NOR2X1_707 ( .A(reset), .B(reg_sh__abc_3798_n72), .Y(reg_sh__abc_3798_n105) );
	NAND2X1 NAND2X1_1102 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n105), .Y(reg_sh__abc_3798_n106) );
	NAND2X1 NAND2X1_1103 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n107) );
	NAND2X1 NAND2X1_1104 ( .A(reg_sh__abc_3798_n107), .B(reg_sh__abc_3798_n106), .Y(reg_sh_value_13__FF_INPUT) );
	NOR2X1 NOR2X1_708 ( .A(reset), .B(reg_sh__abc_3798_n74_1), .Y(reg_sh__abc_3798_n109) );
	NAND2X1 NAND2X1_1105 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n109), .Y(reg_sh__abc_3798_n110) );
	NAND2X1 NAND2X1_1106 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n111) );
	NAND2X1 NAND2X1_1107 ( .A(reg_sh__abc_3798_n111), .B(reg_sh__abc_3798_n110), .Y(reg_sh_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_709 ( .A(reset), .B(reg_sh__abc_3798_n76_1), .Y(reg_sh__abc_3798_n113) );
	NAND2X1 NAND2X1_1108 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n113), .Y(reg_sh__abc_3798_n114) );
	NAND2X1 NAND2X1_1109 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n115) );
	NAND2X1 NAND2X1_1110 ( .A(reg_sh__abc_3798_n115), .B(reg_sh__abc_3798_n114), .Y(reg_sh_value_11__FF_INPUT) );
	NOR2X1 NOR2X1_710 ( .A(reset), .B(reg_sh__abc_3798_n78), .Y(reg_sh__abc_3798_n117) );
	NAND2X1 NAND2X1_1111 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n117), .Y(reg_sh__abc_3798_n118) );
	NAND2X1 NAND2X1_1112 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n119) );
	NAND2X1 NAND2X1_1113 ( .A(reg_sh__abc_3798_n119), .B(reg_sh__abc_3798_n118), .Y(reg_sh_value_10__FF_INPUT) );
	NOR2X1 NOR2X1_711 ( .A(reset), .B(reg_sh__abc_3798_n80_1), .Y(reg_sh__abc_3798_n121) );
	NAND2X1 NAND2X1_1114 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n121), .Y(reg_sh__abc_3798_n122) );
	NAND2X1 NAND2X1_1115 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n123) );
	NAND2X1 NAND2X1_1116 ( .A(reg_sh__abc_3798_n123), .B(reg_sh__abc_3798_n122), .Y(reg_sh_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_712 ( .A(reset), .B(reg_sh__abc_3798_n82_1), .Y(reg_sh__abc_3798_n125) );
	NAND2X1 NAND2X1_1117 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n125), .Y(reg_sh__abc_3798_n126) );
	NAND2X1 NAND2X1_1118 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n127) );
	NAND2X1 NAND2X1_1119 ( .A(reg_sh__abc_3798_n127), .B(reg_sh__abc_3798_n126), .Y(reg_sh_value_8__FF_INPUT) );
	NOR2X1 NOR2X1_713 ( .A(reset), .B(reg_sh__abc_3798_n84_1), .Y(reg_sh__abc_3798_n129) );
	NAND2X1 NAND2X1_1120 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n129), .Y(reg_sh__abc_3798_n130) );
	NAND2X1 NAND2X1_1121 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n131) );
	NAND2X1 NAND2X1_1122 ( .A(reg_sh__abc_3798_n131), .B(reg_sh__abc_3798_n130), .Y(reg_sh_value_7__FF_INPUT) );
	NOR2X1 NOR2X1_714 ( .A(reset), .B(reg_sh__abc_3798_n86), .Y(reg_sh__abc_3798_n133) );
	NAND2X1 NAND2X1_1123 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n133), .Y(reg_sh__abc_3798_n134) );
	NAND2X1 NAND2X1_1124 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n135) );
	NAND2X1 NAND2X1_1125 ( .A(reg_sh__abc_3798_n135), .B(reg_sh__abc_3798_n134), .Y(reg_sh_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_715 ( .A(reset), .B(reg_sh__abc_3798_n88), .Y(reg_sh__abc_3798_n137) );
	NAND2X1 NAND2X1_1126 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n137), .Y(reg_sh__abc_3798_n138) );
	NAND2X1 NAND2X1_1127 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n139) );
	NAND2X1 NAND2X1_1128 ( .A(reg_sh__abc_3798_n139), .B(reg_sh__abc_3798_n138), .Y(reg_sh_value_5__FF_INPUT) );
	NOR2X1 NOR2X1_716 ( .A(reset), .B(reg_sh__abc_3798_n90), .Y(reg_sh__abc_3798_n141) );
	NAND2X1 NAND2X1_1129 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n141), .Y(reg_sh__abc_3798_n142) );
	NAND2X1 NAND2X1_1130 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n143) );
	NAND2X1 NAND2X1_1131 ( .A(reg_sh__abc_3798_n143), .B(reg_sh__abc_3798_n142), .Y(reg_sh_value_4__FF_INPUT) );
	NOR2X1 NOR2X1_717 ( .A(reset), .B(reg_sh__abc_3798_n92), .Y(reg_sh__abc_3798_n145) );
	NAND2X1 NAND2X1_1132 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n145), .Y(reg_sh__abc_3798_n146) );
	NAND2X1 NAND2X1_1133 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n147) );
	NAND2X1 NAND2X1_1134 ( .A(reg_sh__abc_3798_n147), .B(reg_sh__abc_3798_n146), .Y(reg_sh_value_3__FF_INPUT) );
	NOR2X1 NOR2X1_718 ( .A(reset), .B(reg_sh__abc_3798_n94), .Y(reg_sh__abc_3798_n149) );
	NAND2X1 NAND2X1_1135 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n149), .Y(reg_sh__abc_3798_n150) );
	NAND2X1 NAND2X1_1136 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n151) );
	NAND2X1 NAND2X1_1137 ( .A(reg_sh__abc_3798_n151), .B(reg_sh__abc_3798_n150), .Y(reg_sh__abc_3798_n71) );
	NOR2X1 NOR2X1_719 ( .A(reset), .B(reg_sh__abc_3798_n96), .Y(reg_sh__abc_3798_n153) );
	NAND2X1 NAND2X1_1138 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n153), .Y(reg_sh__abc_3798_n154) );
	NAND2X1 NAND2X1_1139 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n155) );
	NAND2X1 NAND2X1_1140 ( .A(reg_sh__abc_3798_n155), .B(reg_sh__abc_3798_n154), .Y(reg_sh__abc_3798_n74) );
	NOR2X1 NOR2X1_720 ( .A(reset), .B(reg_sh__abc_3798_n98), .Y(reg_sh__abc_3798_n157) );
	NAND2X1 NAND2X1_1141 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n157), .Y(reg_sh__abc_3798_n158) );
	NAND2X1 NAND2X1_1142 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n159) );
	NAND2X1 NAND2X1_1143 ( .A(reg_sh__abc_3798_n159), .B(reg_sh__abc_3798_n158), .Y(reg_sh__abc_3798_n77) );
	INVX1 INVX1_288 ( .A(reg_sh_value_15_), .Y(reg_sh__abc_3798_n161) );
	NOR2X1 NOR2X1_721 ( .A(reset), .B(reg_sh__abc_3798_n161), .Y(reg_sh__abc_3798_n162) );
	NAND2X1 NAND2X1_1144 ( .A(reg_sh__abc_3798_n100), .B(reg_sh__abc_3798_n162), .Y(reg_sh__abc_3798_n163) );
	NAND2X1 NAND2X1_1145 ( .A(reset), .B(gnd), .Y(reg_sh__abc_3798_n164) );
	NAND2X1 NAND2X1_1146 ( .A(reg_sh__abc_3798_n164), .B(reg_sh__abc_3798_n163), .Y(reg_sh__abc_3798_n81) );
	NOR2X1 NOR2X1_722 ( .A(reg_sh__abc_3798_n161), .B(reg_sh__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_210 ( .CLK(clk), .D(reg_sh__abc_3798_n77), .Q(reg_sh_value_0_) );
	DFFPOSX1 DFFPOSX1_211 ( .CLK(clk), .D(reg_sh__abc_3798_n74), .Q(reg_sh_value_1_) );
	DFFPOSX1 DFFPOSX1_212 ( .CLK(clk), .D(reg_sh__abc_3798_n71), .Q(reg_sh_value_2_) );
	DFFPOSX1 DFFPOSX1_213 ( .CLK(clk), .D(reg_sh_value_3__FF_INPUT), .Q(reg_sh_value_3_) );
	DFFPOSX1 DFFPOSX1_214 ( .CLK(clk), .D(reg_sh_value_4__FF_INPUT), .Q(reg_sh_value_4_) );
	DFFPOSX1 DFFPOSX1_215 ( .CLK(clk), .D(reg_sh_value_5__FF_INPUT), .Q(reg_sh_value_5_) );
	DFFPOSX1 DFFPOSX1_216 ( .CLK(clk), .D(reg_sh_value_6__FF_INPUT), .Q(reg_sh_value_6_) );
	DFFPOSX1 DFFPOSX1_217 ( .CLK(clk), .D(reg_sh_value_7__FF_INPUT), .Q(reg_sh_value_7_) );
	DFFPOSX1 DFFPOSX1_218 ( .CLK(clk), .D(reg_sh_value_8__FF_INPUT), .Q(reg_sh_value_8_) );
	DFFPOSX1 DFFPOSX1_219 ( .CLK(clk), .D(reg_sh_value_9__FF_INPUT), .Q(reg_sh_value_9_) );
	DFFPOSX1 DFFPOSX1_220 ( .CLK(clk), .D(reg_sh_value_10__FF_INPUT), .Q(reg_sh_value_10_) );
	DFFPOSX1 DFFPOSX1_221 ( .CLK(clk), .D(reg_sh_value_11__FF_INPUT), .Q(reg_sh_value_11_) );
	DFFPOSX1 DFFPOSX1_222 ( .CLK(clk), .D(reg_sh_value_12__FF_INPUT), .Q(reg_sh_value_12_) );
	DFFPOSX1 DFFPOSX1_223 ( .CLK(clk), .D(reg_sh_value_13__FF_INPUT), .Q(reg_sh_value_13_) );
	DFFPOSX1 DFFPOSX1_224 ( .CLK(clk), .D(reg_sh_value_14__FF_INPUT), .Q(reg_sh_value_14_) );
	DFFPOSX1 DFFPOSX1_225 ( .CLK(clk), .D(reg_sh__abc_3798_n81), .Q(reg_sh_value_15_) );
	INVX1 INVX1_289 ( .A(reg_sl_value_14_), .Y(reg_sl__abc_3798_n68_1) );
	INVX1 INVX1_290 ( .A(we), .Y(reg_sl__abc_3798_n69) );
	NAND2X1 NAND2X1_1147 ( .A(addr_sl), .B(reg_sl__abc_3798_n69), .Y(reg_sl__abc_3798_n70_1) );
	NOR2X1 NOR2X1_723 ( .A(reg_sl__abc_3798_n68_1), .B(reg_sl__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_291 ( .A(reg_sl_value_13_), .Y(reg_sl__abc_3798_n72) );
	NOR2X1 NOR2X1_724 ( .A(reg_sl__abc_3798_n72), .B(reg_sl__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_292 ( .A(reg_sl_value_12_), .Y(reg_sl__abc_3798_n74_1) );
	NOR2X1 NOR2X1_725 ( .A(reg_sl__abc_3798_n74_1), .B(reg_sl__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_293 ( .A(reg_sl_value_11_), .Y(reg_sl__abc_3798_n76_1) );
	NOR2X1 NOR2X1_726 ( .A(reg_sl__abc_3798_n76_1), .B(reg_sl__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_294 ( .A(reg_sl_value_10_), .Y(reg_sl__abc_3798_n78) );
	NOR2X1 NOR2X1_727 ( .A(reg_sl__abc_3798_n78), .B(reg_sl__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_295 ( .A(reg_sl_value_9_), .Y(reg_sl__abc_3798_n80_1) );
	NOR2X1 NOR2X1_728 ( .A(reg_sl__abc_3798_n80_1), .B(reg_sl__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_296 ( .A(reg_sl_value_8_), .Y(reg_sl__abc_3798_n82_1) );
	NOR2X1 NOR2X1_729 ( .A(reg_sl__abc_3798_n82_1), .B(reg_sl__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_297 ( .A(reg_sl_value_7_), .Y(reg_sl__abc_3798_n84_1) );
	NOR2X1 NOR2X1_730 ( .A(reg_sl__abc_3798_n84_1), .B(reg_sl__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_298 ( .A(reg_sl_value_6_), .Y(reg_sl__abc_3798_n86) );
	NOR2X1 NOR2X1_731 ( .A(reg_sl__abc_3798_n86), .B(reg_sl__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_299 ( .A(reg_sl_value_5_), .Y(reg_sl__abc_3798_n88) );
	NOR2X1 NOR2X1_732 ( .A(reg_sl__abc_3798_n88), .B(reg_sl__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_300 ( .A(reg_sl_value_4_), .Y(reg_sl__abc_3798_n90) );
	NOR2X1 NOR2X1_733 ( .A(reg_sl__abc_3798_n90), .B(reg_sl__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_301 ( .A(reg_sl_value_3_), .Y(reg_sl__abc_3798_n92) );
	NOR2X1 NOR2X1_734 ( .A(reg_sl__abc_3798_n92), .B(reg_sl__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_302 ( .A(reg_sl_value_2_), .Y(reg_sl__abc_3798_n94) );
	NOR2X1 NOR2X1_735 ( .A(reg_sl__abc_3798_n94), .B(reg_sl__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_303 ( .A(reg_sl_value_1_), .Y(reg_sl__abc_3798_n96) );
	NOR2X1 NOR2X1_736 ( .A(reg_sl__abc_3798_n96), .B(reg_sl__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_304 ( .A(reg_sl_value_0_), .Y(reg_sl__abc_3798_n98) );
	NOR2X1 NOR2X1_737 ( .A(reg_sl__abc_3798_n98), .B(reg_sl__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1148 ( .A(we), .B(addr_sl), .Y(reg_sl__abc_3798_n100) );
	NOR2X1 NOR2X1_738 ( .A(reset), .B(reg_sl__abc_3798_n68_1), .Y(reg_sl__abc_3798_n101) );
	NAND2X1 NAND2X1_1149 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n101), .Y(reg_sl__abc_3798_n102) );
	NAND2X1 NAND2X1_1150 ( .A(gnd), .B(reset), .Y(reg_sl__abc_3798_n103) );
	NAND2X1 NAND2X1_1151 ( .A(reg_sl__abc_3798_n103), .B(reg_sl__abc_3798_n102), .Y(reg_sl__abc_3798_n35) );
	NOR2X1 NOR2X1_739 ( .A(reset), .B(reg_sl__abc_3798_n72), .Y(reg_sl__abc_3798_n105) );
	NAND2X1 NAND2X1_1152 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n105), .Y(reg_sl__abc_3798_n106) );
	NAND2X1 NAND2X1_1153 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n107) );
	NAND2X1 NAND2X1_1154 ( .A(reg_sl__abc_3798_n107), .B(reg_sl__abc_3798_n106), .Y(reg_sl__abc_3798_n38) );
	NOR2X1 NOR2X1_740 ( .A(reset), .B(reg_sl__abc_3798_n74_1), .Y(reg_sl__abc_3798_n109) );
	NAND2X1 NAND2X1_1155 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n109), .Y(reg_sl__abc_3798_n110) );
	NAND2X1 NAND2X1_1156 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n111) );
	NAND2X1 NAND2X1_1157 ( .A(reg_sl__abc_3798_n111), .B(reg_sl__abc_3798_n110), .Y(reg_sl__abc_3798_n41) );
	NOR2X1 NOR2X1_741 ( .A(reset), .B(reg_sl__abc_3798_n76_1), .Y(reg_sl__abc_3798_n113) );
	NAND2X1 NAND2X1_1158 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n113), .Y(reg_sl__abc_3798_n114) );
	NAND2X1 NAND2X1_1159 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n115) );
	NAND2X1 NAND2X1_1160 ( .A(reg_sl__abc_3798_n115), .B(reg_sl__abc_3798_n114), .Y(reg_sl__abc_3798_n44) );
	NOR2X1 NOR2X1_742 ( .A(reset), .B(reg_sl__abc_3798_n78), .Y(reg_sl__abc_3798_n117) );
	NAND2X1 NAND2X1_1161 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n117), .Y(reg_sl__abc_3798_n118) );
	NAND2X1 NAND2X1_1162 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n119) );
	NAND2X1 NAND2X1_1163 ( .A(reg_sl__abc_3798_n119), .B(reg_sl__abc_3798_n118), .Y(reg_sl__abc_3798_n47) );
	NOR2X1 NOR2X1_743 ( .A(reset), .B(reg_sl__abc_3798_n80_1), .Y(reg_sl__abc_3798_n121) );
	NAND2X1 NAND2X1_1164 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n121), .Y(reg_sl__abc_3798_n122) );
	NAND2X1 NAND2X1_1165 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n123) );
	NAND2X1 NAND2X1_1166 ( .A(reg_sl__abc_3798_n123), .B(reg_sl__abc_3798_n122), .Y(reg_sl__abc_3798_n50) );
	NOR2X1 NOR2X1_744 ( .A(reset), .B(reg_sl__abc_3798_n82_1), .Y(reg_sl__abc_3798_n125) );
	NAND2X1 NAND2X1_1167 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n125), .Y(reg_sl__abc_3798_n126) );
	NAND2X1 NAND2X1_1168 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n127) );
	NAND2X1 NAND2X1_1169 ( .A(reg_sl__abc_3798_n127), .B(reg_sl__abc_3798_n126), .Y(reg_sl__abc_3798_n53) );
	NOR2X1 NOR2X1_745 ( .A(reset), .B(reg_sl__abc_3798_n84_1), .Y(reg_sl__abc_3798_n129) );
	NAND2X1 NAND2X1_1170 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n129), .Y(reg_sl__abc_3798_n130) );
	NAND2X1 NAND2X1_1171 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n131) );
	NAND2X1 NAND2X1_1172 ( .A(reg_sl__abc_3798_n131), .B(reg_sl__abc_3798_n130), .Y(reg_sl__abc_3798_n56) );
	NOR2X1 NOR2X1_746 ( .A(reset), .B(reg_sl__abc_3798_n86), .Y(reg_sl__abc_3798_n133) );
	NAND2X1 NAND2X1_1173 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n133), .Y(reg_sl__abc_3798_n134) );
	NAND2X1 NAND2X1_1174 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n135) );
	NAND2X1 NAND2X1_1175 ( .A(reg_sl__abc_3798_n135), .B(reg_sl__abc_3798_n134), .Y(reg_sl__abc_3798_n59) );
	NOR2X1 NOR2X1_747 ( .A(reset), .B(reg_sl__abc_3798_n88), .Y(reg_sl__abc_3798_n137) );
	NAND2X1 NAND2X1_1176 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n137), .Y(reg_sl__abc_3798_n138) );
	NAND2X1 NAND2X1_1177 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n139) );
	NAND2X1 NAND2X1_1178 ( .A(reg_sl__abc_3798_n139), .B(reg_sl__abc_3798_n138), .Y(reg_sl__abc_3798_n62) );
	NOR2X1 NOR2X1_748 ( .A(reset), .B(reg_sl__abc_3798_n90), .Y(reg_sl__abc_3798_n141) );
	NAND2X1 NAND2X1_1179 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n141), .Y(reg_sl__abc_3798_n142) );
	NAND2X1 NAND2X1_1180 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n143) );
	NAND2X1 NAND2X1_1181 ( .A(reg_sl__abc_3798_n143), .B(reg_sl__abc_3798_n142), .Y(reg_sl__abc_3798_n65) );
	NOR2X1 NOR2X1_749 ( .A(reset), .B(reg_sl__abc_3798_n92), .Y(reg_sl__abc_3798_n145) );
	NAND2X1 NAND2X1_1182 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n145), .Y(reg_sl__abc_3798_n146) );
	NAND2X1 NAND2X1_1183 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n147) );
	NAND2X1 NAND2X1_1184 ( .A(reg_sl__abc_3798_n147), .B(reg_sl__abc_3798_n146), .Y(reg_sl__abc_3798_n68) );
	NOR2X1 NOR2X1_750 ( .A(reset), .B(reg_sl__abc_3798_n94), .Y(reg_sl__abc_3798_n149) );
	NAND2X1 NAND2X1_1185 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n149), .Y(reg_sl__abc_3798_n150) );
	NAND2X1 NAND2X1_1186 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n151) );
	NAND2X1 NAND2X1_1187 ( .A(reg_sl__abc_3798_n151), .B(reg_sl__abc_3798_n150), .Y(reg_sl__abc_3798_n71) );
	NOR2X1 NOR2X1_751 ( .A(reset), .B(reg_sl__abc_3798_n96), .Y(reg_sl__abc_3798_n153) );
	NAND2X1 NAND2X1_1188 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n153), .Y(reg_sl__abc_3798_n154) );
	NAND2X1 NAND2X1_1189 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n155) );
	NAND2X1 NAND2X1_1190 ( .A(reg_sl__abc_3798_n155), .B(reg_sl__abc_3798_n154), .Y(reg_sl__abc_3798_n74) );
	NOR2X1 NOR2X1_752 ( .A(reset), .B(reg_sl__abc_3798_n98), .Y(reg_sl__abc_3798_n157) );
	NAND2X1 NAND2X1_1191 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n157), .Y(reg_sl__abc_3798_n158) );
	NAND2X1 NAND2X1_1192 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n159) );
	NAND2X1 NAND2X1_1193 ( .A(reg_sl__abc_3798_n159), .B(reg_sl__abc_3798_n158), .Y(reg_sl__abc_3798_n77) );
	INVX1 INVX1_305 ( .A(reg_sl_value_15_), .Y(reg_sl__abc_3798_n161) );
	NOR2X1 NOR2X1_753 ( .A(reset), .B(reg_sl__abc_3798_n161), .Y(reg_sl__abc_3798_n162) );
	NAND2X1 NAND2X1_1194 ( .A(reg_sl__abc_3798_n100), .B(reg_sl__abc_3798_n162), .Y(reg_sl__abc_3798_n163) );
	NAND2X1 NAND2X1_1195 ( .A(reset), .B(gnd), .Y(reg_sl__abc_3798_n164) );
	NAND2X1 NAND2X1_1196 ( .A(reg_sl__abc_3798_n164), .B(reg_sl__abc_3798_n163), .Y(reg_sl__abc_3798_n81) );
	NOR2X1 NOR2X1_754 ( .A(reg_sl__abc_3798_n161), .B(reg_sl__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_226 ( .CLK(clk), .D(reg_sl__abc_3798_n77), .Q(reg_sl_value_0_) );
	DFFPOSX1 DFFPOSX1_227 ( .CLK(clk), .D(reg_sl__abc_3798_n74), .Q(reg_sl_value_1_) );
	DFFPOSX1 DFFPOSX1_228 ( .CLK(clk), .D(reg_sl__abc_3798_n71), .Q(reg_sl_value_2_) );
	DFFPOSX1 DFFPOSX1_229 ( .CLK(clk), .D(reg_sl__abc_3798_n68), .Q(reg_sl_value_3_) );
	DFFPOSX1 DFFPOSX1_230 ( .CLK(clk), .D(reg_sl__abc_3798_n65), .Q(reg_sl_value_4_) );
	DFFPOSX1 DFFPOSX1_231 ( .CLK(clk), .D(reg_sl__abc_3798_n62), .Q(reg_sl_value_5_) );
	DFFPOSX1 DFFPOSX1_232 ( .CLK(clk), .D(reg_sl__abc_3798_n59), .Q(reg_sl_value_6_) );
	DFFPOSX1 DFFPOSX1_233 ( .CLK(clk), .D(reg_sl__abc_3798_n56), .Q(reg_sl_value_7_) );
	DFFPOSX1 DFFPOSX1_234 ( .CLK(clk), .D(reg_sl__abc_3798_n53), .Q(reg_sl_value_8_) );
	DFFPOSX1 DFFPOSX1_235 ( .CLK(clk), .D(reg_sl__abc_3798_n50), .Q(reg_sl_value_9_) );
	DFFPOSX1 DFFPOSX1_236 ( .CLK(clk), .D(reg_sl__abc_3798_n47), .Q(reg_sl_value_10_) );
	DFFPOSX1 DFFPOSX1_237 ( .CLK(clk), .D(reg_sl__abc_3798_n44), .Q(reg_sl_value_11_) );
	DFFPOSX1 DFFPOSX1_238 ( .CLK(clk), .D(reg_sl__abc_3798_n41), .Q(reg_sl_value_12_) );
	DFFPOSX1 DFFPOSX1_239 ( .CLK(clk), .D(reg_sl__abc_3798_n38), .Q(reg_sl_value_13_) );
	DFFPOSX1 DFFPOSX1_240 ( .CLK(clk), .D(reg_sl__abc_3798_n35), .Q(reg_sl_value_14_) );
	DFFPOSX1 DFFPOSX1_241 ( .CLK(clk), .D(reg_sl__abc_3798_n81), .Q(reg_sl_value_15_) );
	INVX1 INVX1_306 ( .A(reg_vb_value_14_), .Y(reg_vb__abc_3798_n68_1) );
	INVX1 INVX1_307 ( .A(we), .Y(reg_vb__abc_3798_n69) );
	NAND2X1 NAND2X1_1197 ( .A(addr_vb), .B(reg_vb__abc_3798_n69), .Y(reg_vb__abc_3798_n70_1) );
	NOR2X1 NOR2X1_755 ( .A(reg_vb__abc_3798_n68_1), .B(reg_vb__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_308 ( .A(reg_vb_value_13_), .Y(reg_vb__abc_3798_n72) );
	NOR2X1 NOR2X1_756 ( .A(reg_vb__abc_3798_n72), .B(reg_vb__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_309 ( .A(reg_vb_value_12_), .Y(reg_vb__abc_3798_n74_1) );
	NOR2X1 NOR2X1_757 ( .A(reg_vb__abc_3798_n74_1), .B(reg_vb__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_310 ( .A(reg_vb_value_11_), .Y(reg_vb__abc_3798_n76_1) );
	NOR2X1 NOR2X1_758 ( .A(reg_vb__abc_3798_n76_1), .B(reg_vb__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_311 ( .A(reg_vb_value_10_), .Y(reg_vb__abc_3798_n78) );
	NOR2X1 NOR2X1_759 ( .A(reg_vb__abc_3798_n78), .B(reg_vb__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_312 ( .A(reg_vb_value_9_), .Y(reg_vb__abc_3798_n80_1) );
	NOR2X1 NOR2X1_760 ( .A(reg_vb__abc_3798_n80_1), .B(reg_vb__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_313 ( .A(reg_vb_value_8_), .Y(reg_vb__abc_3798_n82_1) );
	NOR2X1 NOR2X1_761 ( .A(reg_vb__abc_3798_n82_1), .B(reg_vb__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_314 ( .A(reg_vb_value_7_), .Y(reg_vb__abc_3798_n84_1) );
	NOR2X1 NOR2X1_762 ( .A(reg_vb__abc_3798_n84_1), .B(reg_vb__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_315 ( .A(reg_vb_value_6_), .Y(reg_vb__abc_3798_n86) );
	NOR2X1 NOR2X1_763 ( .A(reg_vb__abc_3798_n86), .B(reg_vb__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_316 ( .A(reg_vb_value_5_), .Y(reg_vb__abc_3798_n88) );
	NOR2X1 NOR2X1_764 ( .A(reg_vb__abc_3798_n88), .B(reg_vb__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_317 ( .A(reg_vb_value_4_), .Y(reg_vb__abc_3798_n90) );
	NOR2X1 NOR2X1_765 ( .A(reg_vb__abc_3798_n90), .B(reg_vb__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_318 ( .A(reg_vb_value_3_), .Y(reg_vb__abc_3798_n92) );
	NOR2X1 NOR2X1_766 ( .A(reg_vb__abc_3798_n92), .B(reg_vb__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_319 ( .A(reg_vb_value_2_), .Y(reg_vb__abc_3798_n94) );
	NOR2X1 NOR2X1_767 ( .A(reg_vb__abc_3798_n94), .B(reg_vb__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_320 ( .A(reg_vb_value_1_), .Y(reg_vb__abc_3798_n96) );
	NOR2X1 NOR2X1_768 ( .A(reg_vb__abc_3798_n96), .B(reg_vb__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_321 ( .A(reg_vb_value_0_), .Y(reg_vb__abc_3798_n98) );
	NOR2X1 NOR2X1_769 ( .A(reg_vb__abc_3798_n98), .B(reg_vb__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1198 ( .A(we), .B(addr_vb), .Y(reg_vb__abc_3798_n100) );
	NOR2X1 NOR2X1_770 ( .A(reset), .B(reg_vb__abc_3798_n68_1), .Y(reg_vb__abc_3798_n101) );
	NAND2X1 NAND2X1_1199 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n101), .Y(reg_vb__abc_3798_n102) );
	NAND2X1 NAND2X1_1200 ( .A(gnd), .B(reset), .Y(reg_vb__abc_3798_n103) );
	NAND2X1 NAND2X1_1201 ( .A(reg_vb__abc_3798_n103), .B(reg_vb__abc_3798_n102), .Y(reg_vb__abc_3798_n35) );
	NOR2X1 NOR2X1_771 ( .A(reset), .B(reg_vb__abc_3798_n72), .Y(reg_vb__abc_3798_n105) );
	NAND2X1 NAND2X1_1202 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n105), .Y(reg_vb__abc_3798_n106) );
	NAND2X1 NAND2X1_1203 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n107) );
	NAND2X1 NAND2X1_1204 ( .A(reg_vb__abc_3798_n107), .B(reg_vb__abc_3798_n106), .Y(reg_vb__abc_3798_n38) );
	NOR2X1 NOR2X1_772 ( .A(reset), .B(reg_vb__abc_3798_n74_1), .Y(reg_vb__abc_3798_n109) );
	NAND2X1 NAND2X1_1205 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n109), .Y(reg_vb__abc_3798_n110) );
	NAND2X1 NAND2X1_1206 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n111) );
	NAND2X1 NAND2X1_1207 ( .A(reg_vb__abc_3798_n111), .B(reg_vb__abc_3798_n110), .Y(reg_vb__abc_3798_n41) );
	NOR2X1 NOR2X1_773 ( .A(reset), .B(reg_vb__abc_3798_n76_1), .Y(reg_vb__abc_3798_n113) );
	NAND2X1 NAND2X1_1208 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n113), .Y(reg_vb__abc_3798_n114) );
	NAND2X1 NAND2X1_1209 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n115) );
	NAND2X1 NAND2X1_1210 ( .A(reg_vb__abc_3798_n115), .B(reg_vb__abc_3798_n114), .Y(reg_vb__abc_3798_n44) );
	NOR2X1 NOR2X1_774 ( .A(reset), .B(reg_vb__abc_3798_n78), .Y(reg_vb__abc_3798_n117) );
	NAND2X1 NAND2X1_1211 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n117), .Y(reg_vb__abc_3798_n118) );
	NAND2X1 NAND2X1_1212 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n119) );
	NAND2X1 NAND2X1_1213 ( .A(reg_vb__abc_3798_n119), .B(reg_vb__abc_3798_n118), .Y(reg_vb__abc_3798_n47) );
	NOR2X1 NOR2X1_775 ( .A(reset), .B(reg_vb__abc_3798_n80_1), .Y(reg_vb__abc_3798_n121) );
	NAND2X1 NAND2X1_1214 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n121), .Y(reg_vb__abc_3798_n122) );
	NAND2X1 NAND2X1_1215 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n123) );
	NAND2X1 NAND2X1_1216 ( .A(reg_vb__abc_3798_n123), .B(reg_vb__abc_3798_n122), .Y(reg_vb__abc_3798_n50) );
	NOR2X1 NOR2X1_776 ( .A(reset), .B(reg_vb__abc_3798_n82_1), .Y(reg_vb__abc_3798_n125) );
	NAND2X1 NAND2X1_1217 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n125), .Y(reg_vb__abc_3798_n126) );
	NAND2X1 NAND2X1_1218 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n127) );
	NAND2X1 NAND2X1_1219 ( .A(reg_vb__abc_3798_n127), .B(reg_vb__abc_3798_n126), .Y(reg_vb__abc_3798_n53) );
	NOR2X1 NOR2X1_777 ( .A(reset), .B(reg_vb__abc_3798_n84_1), .Y(reg_vb__abc_3798_n129) );
	NAND2X1 NAND2X1_1220 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n129), .Y(reg_vb__abc_3798_n130) );
	NAND2X1 NAND2X1_1221 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n131) );
	NAND2X1 NAND2X1_1222 ( .A(reg_vb__abc_3798_n131), .B(reg_vb__abc_3798_n130), .Y(reg_vb__abc_3798_n56) );
	NOR2X1 NOR2X1_778 ( .A(reset), .B(reg_vb__abc_3798_n86), .Y(reg_vb__abc_3798_n133) );
	NAND2X1 NAND2X1_1223 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n133), .Y(reg_vb__abc_3798_n134) );
	NAND2X1 NAND2X1_1224 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n135) );
	NAND2X1 NAND2X1_1225 ( .A(reg_vb__abc_3798_n135), .B(reg_vb__abc_3798_n134), .Y(reg_vb__abc_3798_n59) );
	NOR2X1 NOR2X1_779 ( .A(reset), .B(reg_vb__abc_3798_n88), .Y(reg_vb__abc_3798_n137) );
	NAND2X1 NAND2X1_1226 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n137), .Y(reg_vb__abc_3798_n138) );
	NAND2X1 NAND2X1_1227 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n139) );
	NAND2X1 NAND2X1_1228 ( .A(reg_vb__abc_3798_n139), .B(reg_vb__abc_3798_n138), .Y(reg_vb__abc_3798_n62) );
	NOR2X1 NOR2X1_780 ( .A(reset), .B(reg_vb__abc_3798_n90), .Y(reg_vb__abc_3798_n141) );
	NAND2X1 NAND2X1_1229 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n141), .Y(reg_vb__abc_3798_n142) );
	NAND2X1 NAND2X1_1230 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n143) );
	NAND2X1 NAND2X1_1231 ( .A(reg_vb__abc_3798_n143), .B(reg_vb__abc_3798_n142), .Y(reg_vb__abc_3798_n65) );
	NOR2X1 NOR2X1_781 ( .A(reset), .B(reg_vb__abc_3798_n92), .Y(reg_vb__abc_3798_n145) );
	NAND2X1 NAND2X1_1232 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n145), .Y(reg_vb__abc_3798_n146) );
	NAND2X1 NAND2X1_1233 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n147) );
	NAND2X1 NAND2X1_1234 ( .A(reg_vb__abc_3798_n147), .B(reg_vb__abc_3798_n146), .Y(reg_vb__abc_3798_n68) );
	NOR2X1 NOR2X1_782 ( .A(reset), .B(reg_vb__abc_3798_n94), .Y(reg_vb__abc_3798_n149) );
	NAND2X1 NAND2X1_1235 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n149), .Y(reg_vb__abc_3798_n150) );
	NAND2X1 NAND2X1_1236 ( .A(reset), .B(vdd), .Y(reg_vb__abc_3798_n151) );
	NAND2X1 NAND2X1_1237 ( .A(reg_vb__abc_3798_n151), .B(reg_vb__abc_3798_n150), .Y(reg_vb__abc_3798_n71) );
	NOR2X1 NOR2X1_783 ( .A(reset), .B(reg_vb__abc_3798_n96), .Y(reg_vb__abc_3798_n153) );
	NAND2X1 NAND2X1_1238 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n153), .Y(reg_vb__abc_3798_n154) );
	NAND2X1 NAND2X1_1239 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n155) );
	NAND2X1 NAND2X1_1240 ( .A(reg_vb__abc_3798_n155), .B(reg_vb__abc_3798_n154), .Y(reg_vb__abc_3798_n74) );
	NOR2X1 NOR2X1_784 ( .A(reset), .B(reg_vb__abc_3798_n98), .Y(reg_vb__abc_3798_n157) );
	NAND2X1 NAND2X1_1241 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n157), .Y(reg_vb__abc_3798_n158) );
	NAND2X1 NAND2X1_1242 ( .A(reset), .B(vdd), .Y(reg_vb__abc_3798_n159) );
	NAND2X1 NAND2X1_1243 ( .A(reg_vb__abc_3798_n159), .B(reg_vb__abc_3798_n158), .Y(reg_vb__abc_3798_n77) );
	INVX1 INVX1_322 ( .A(reg_vb_value_15_), .Y(reg_vb__abc_3798_n161) );
	NOR2X1 NOR2X1_785 ( .A(reset), .B(reg_vb__abc_3798_n161), .Y(reg_vb__abc_3798_n162) );
	NAND2X1 NAND2X1_1244 ( .A(reg_vb__abc_3798_n100), .B(reg_vb__abc_3798_n162), .Y(reg_vb__abc_3798_n163) );
	NAND2X1 NAND2X1_1245 ( .A(reset), .B(gnd), .Y(reg_vb__abc_3798_n164) );
	NAND2X1 NAND2X1_1246 ( .A(reg_vb__abc_3798_n164), .B(reg_vb__abc_3798_n163), .Y(reg_vb__abc_3798_n81) );
	NOR2X1 NOR2X1_786 ( .A(reg_vb__abc_3798_n161), .B(reg_vb__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_242 ( .CLK(clk), .D(reg_vb__abc_3798_n77), .Q(reg_vb_value_0_) );
	DFFPOSX1 DFFPOSX1_243 ( .CLK(clk), .D(reg_vb__abc_3798_n74), .Q(reg_vb_value_1_) );
	DFFPOSX1 DFFPOSX1_244 ( .CLK(clk), .D(reg_vb__abc_3798_n71), .Q(reg_vb_value_2_) );
	DFFPOSX1 DFFPOSX1_245 ( .CLK(clk), .D(reg_vb__abc_3798_n68), .Q(reg_vb_value_3_) );
	DFFPOSX1 DFFPOSX1_246 ( .CLK(clk), .D(reg_vb__abc_3798_n65), .Q(reg_vb_value_4_) );
	DFFPOSX1 DFFPOSX1_247 ( .CLK(clk), .D(reg_vb__abc_3798_n62), .Q(reg_vb_value_5_) );
	DFFPOSX1 DFFPOSX1_248 ( .CLK(clk), .D(reg_vb__abc_3798_n59), .Q(reg_vb_value_6_) );
	DFFPOSX1 DFFPOSX1_249 ( .CLK(clk), .D(reg_vb__abc_3798_n56), .Q(reg_vb_value_7_) );
	DFFPOSX1 DFFPOSX1_250 ( .CLK(clk), .D(reg_vb__abc_3798_n53), .Q(reg_vb_value_8_) );
	DFFPOSX1 DFFPOSX1_251 ( .CLK(clk), .D(reg_vb__abc_3798_n50), .Q(reg_vb_value_9_) );
	DFFPOSX1 DFFPOSX1_252 ( .CLK(clk), .D(reg_vb__abc_3798_n47), .Q(reg_vb_value_10_) );
	DFFPOSX1 DFFPOSX1_253 ( .CLK(clk), .D(reg_vb__abc_3798_n44), .Q(reg_vb_value_11_) );
	DFFPOSX1 DFFPOSX1_254 ( .CLK(clk), .D(reg_vb__abc_3798_n41), .Q(reg_vb_value_12_) );
	DFFPOSX1 DFFPOSX1_255 ( .CLK(clk), .D(reg_vb__abc_3798_n38), .Q(reg_vb_value_13_) );
	DFFPOSX1 DFFPOSX1_256 ( .CLK(clk), .D(reg_vb__abc_3798_n35), .Q(reg_vb_value_14_) );
	DFFPOSX1 DFFPOSX1_257 ( .CLK(clk), .D(reg_vb__abc_3798_n81), .Q(reg_vb_value_15_) );
	INVX1 INVX1_323 ( .A(reg_ve_value_14_), .Y(reg_ve__abc_3798_n68_1) );
	INVX1 INVX1_324 ( .A(we), .Y(reg_ve__abc_3798_n69) );
	NAND2X1 NAND2X1_1247 ( .A(addr_ve), .B(reg_ve__abc_3798_n69), .Y(reg_ve__abc_3798_n70_1) );
	NOR2X1 NOR2X1_787 ( .A(reg_ve__abc_3798_n68_1), .B(reg_ve__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_325 ( .A(reg_ve_value_13_), .Y(reg_ve__abc_3798_n72) );
	NOR2X1 NOR2X1_788 ( .A(reg_ve__abc_3798_n72), .B(reg_ve__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_326 ( .A(reg_ve_value_12_), .Y(reg_ve__abc_3798_n74_1) );
	NOR2X1 NOR2X1_789 ( .A(reg_ve__abc_3798_n74_1), .B(reg_ve__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_327 ( .A(reg_ve_value_11_), .Y(reg_ve__abc_3798_n76_1) );
	NOR2X1 NOR2X1_790 ( .A(reg_ve__abc_3798_n76_1), .B(reg_ve__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_328 ( .A(reg_ve_value_10_), .Y(reg_ve__abc_3798_n78) );
	NOR2X1 NOR2X1_791 ( .A(reg_ve__abc_3798_n78), .B(reg_ve__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_329 ( .A(reg_ve_value_9_), .Y(reg_ve__abc_3798_n80_1) );
	NOR2X1 NOR2X1_792 ( .A(reg_ve__abc_3798_n80_1), .B(reg_ve__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_330 ( .A(reg_ve_value_8_), .Y(reg_ve__abc_3798_n82_1) );
	NOR2X1 NOR2X1_793 ( .A(reg_ve__abc_3798_n82_1), .B(reg_ve__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_331 ( .A(reg_ve_value_7_), .Y(reg_ve__abc_3798_n84_1) );
	NOR2X1 NOR2X1_794 ( .A(reg_ve__abc_3798_n84_1), .B(reg_ve__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_332 ( .A(reg_ve_value_6_), .Y(reg_ve__abc_3798_n86) );
	NOR2X1 NOR2X1_795 ( .A(reg_ve__abc_3798_n86), .B(reg_ve__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_333 ( .A(reg_ve_value_5_), .Y(reg_ve__abc_3798_n88) );
	NOR2X1 NOR2X1_796 ( .A(reg_ve__abc_3798_n88), .B(reg_ve__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_334 ( .A(reg_ve_value_4_), .Y(reg_ve__abc_3798_n90) );
	NOR2X1 NOR2X1_797 ( .A(reg_ve__abc_3798_n90), .B(reg_ve__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_335 ( .A(reg_ve_value_3_), .Y(reg_ve__abc_3798_n92) );
	NOR2X1 NOR2X1_798 ( .A(reg_ve__abc_3798_n92), .B(reg_ve__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_336 ( .A(reg_ve_value_2_), .Y(reg_ve__abc_3798_n94) );
	NOR2X1 NOR2X1_799 ( .A(reg_ve__abc_3798_n94), .B(reg_ve__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_337 ( .A(reg_ve_value_1_), .Y(reg_ve__abc_3798_n96) );
	NOR2X1 NOR2X1_800 ( .A(reg_ve__abc_3798_n96), .B(reg_ve__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_338 ( .A(reg_ve_value_0_), .Y(reg_ve__abc_3798_n98) );
	NOR2X1 NOR2X1_801 ( .A(reg_ve__abc_3798_n98), .B(reg_ve__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1248 ( .A(we), .B(addr_ve), .Y(reg_ve__abc_3798_n100) );
	NOR2X1 NOR2X1_802 ( .A(reset), .B(reg_ve__abc_3798_n68_1), .Y(reg_ve__abc_3798_n101) );
	NAND2X1 NAND2X1_1249 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n101), .Y(reg_ve__abc_3798_n102) );
	NAND2X1 NAND2X1_1250 ( .A(gnd), .B(reset), .Y(reg_ve__abc_3798_n103) );
	NAND2X1 NAND2X1_1251 ( .A(reg_ve__abc_3798_n103), .B(reg_ve__abc_3798_n102), .Y(reg_ve__abc_3798_n35) );
	NOR2X1 NOR2X1_803 ( .A(reset), .B(reg_ve__abc_3798_n72), .Y(reg_ve__abc_3798_n105) );
	NAND2X1 NAND2X1_1252 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n105), .Y(reg_ve__abc_3798_n106) );
	NAND2X1 NAND2X1_1253 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n107) );
	NAND2X1 NAND2X1_1254 ( .A(reg_ve__abc_3798_n107), .B(reg_ve__abc_3798_n106), .Y(reg_ve_value_13__FF_INPUT) );
	NOR2X1 NOR2X1_804 ( .A(reset), .B(reg_ve__abc_3798_n74_1), .Y(reg_ve__abc_3798_n109) );
	NAND2X1 NAND2X1_1255 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n109), .Y(reg_ve__abc_3798_n110) );
	NAND2X1 NAND2X1_1256 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n111) );
	NAND2X1 NAND2X1_1257 ( .A(reg_ve__abc_3798_n111), .B(reg_ve__abc_3798_n110), .Y(reg_ve_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_805 ( .A(reset), .B(reg_ve__abc_3798_n76_1), .Y(reg_ve__abc_3798_n113) );
	NAND2X1 NAND2X1_1258 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n113), .Y(reg_ve__abc_3798_n114) );
	NAND2X1 NAND2X1_1259 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n115) );
	NAND2X1 NAND2X1_1260 ( .A(reg_ve__abc_3798_n115), .B(reg_ve__abc_3798_n114), .Y(reg_ve__abc_3798_n44) );
	NOR2X1 NOR2X1_806 ( .A(reset), .B(reg_ve__abc_3798_n78), .Y(reg_ve__abc_3798_n117) );
	NAND2X1 NAND2X1_1261 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n117), .Y(reg_ve__abc_3798_n118) );
	NAND2X1 NAND2X1_1262 ( .A(reset), .B(vdd), .Y(reg_ve__abc_3798_n119) );
	NAND2X1 NAND2X1_1263 ( .A(reg_ve__abc_3798_n119), .B(reg_ve__abc_3798_n118), .Y(reg_ve__abc_3798_n47) );
	NOR2X1 NOR2X1_807 ( .A(reset), .B(reg_ve__abc_3798_n80_1), .Y(reg_ve__abc_3798_n121) );
	NAND2X1 NAND2X1_1264 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n121), .Y(reg_ve__abc_3798_n122) );
	NAND2X1 NAND2X1_1265 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n123) );
	NAND2X1 NAND2X1_1266 ( .A(reg_ve__abc_3798_n123), .B(reg_ve__abc_3798_n122), .Y(reg_ve_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_808 ( .A(reset), .B(reg_ve__abc_3798_n82_1), .Y(reg_ve__abc_3798_n125) );
	NAND2X1 NAND2X1_1267 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n125), .Y(reg_ve__abc_3798_n126) );
	NAND2X1 NAND2X1_1268 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n127) );
	NAND2X1 NAND2X1_1269 ( .A(reg_ve__abc_3798_n127), .B(reg_ve__abc_3798_n126), .Y(reg_ve__abc_3798_n53) );
	NOR2X1 NOR2X1_809 ( .A(reset), .B(reg_ve__abc_3798_n84_1), .Y(reg_ve__abc_3798_n129) );
	NAND2X1 NAND2X1_1270 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n129), .Y(reg_ve__abc_3798_n130) );
	NAND2X1 NAND2X1_1271 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n131) );
	NAND2X1 NAND2X1_1272 ( .A(reg_ve__abc_3798_n131), .B(reg_ve__abc_3798_n130), .Y(reg_ve__abc_3798_n56) );
	NOR2X1 NOR2X1_810 ( .A(reset), .B(reg_ve__abc_3798_n86), .Y(reg_ve__abc_3798_n133) );
	NAND2X1 NAND2X1_1273 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n133), .Y(reg_ve__abc_3798_n134) );
	NAND2X1 NAND2X1_1274 ( .A(reset), .B(vdd), .Y(reg_ve__abc_3798_n135) );
	NAND2X1 NAND2X1_1275 ( .A(reg_ve__abc_3798_n135), .B(reg_ve__abc_3798_n134), .Y(reg_ve_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_811 ( .A(reset), .B(reg_ve__abc_3798_n88), .Y(reg_ve__abc_3798_n137) );
	NAND2X1 NAND2X1_1276 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n137), .Y(reg_ve__abc_3798_n138) );
	NAND2X1 NAND2X1_1277 ( .A(reset), .B(vdd), .Y(reg_ve__abc_3798_n139) );
	NAND2X1 NAND2X1_1278 ( .A(reg_ve__abc_3798_n139), .B(reg_ve__abc_3798_n138), .Y(reg_ve_value_5__FF_INPUT) );
	NOR2X1 NOR2X1_812 ( .A(reset), .B(reg_ve__abc_3798_n90), .Y(reg_ve__abc_3798_n141) );
	NAND2X1 NAND2X1_1279 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n141), .Y(reg_ve__abc_3798_n142) );
	NAND2X1 NAND2X1_1280 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n143) );
	NAND2X1 NAND2X1_1281 ( .A(reg_ve__abc_3798_n143), .B(reg_ve__abc_3798_n142), .Y(reg_ve__abc_3798_n65) );
	NOR2X1 NOR2X1_813 ( .A(reset), .B(reg_ve__abc_3798_n92), .Y(reg_ve__abc_3798_n145) );
	NAND2X1 NAND2X1_1282 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n145), .Y(reg_ve__abc_3798_n146) );
	NAND2X1 NAND2X1_1283 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n147) );
	NAND2X1 NAND2X1_1284 ( .A(reg_ve__abc_3798_n147), .B(reg_ve__abc_3798_n146), .Y(reg_ve_value_3__FF_INPUT) );
	NOR2X1 NOR2X1_814 ( .A(reset), .B(reg_ve__abc_3798_n94), .Y(reg_ve__abc_3798_n149) );
	NAND2X1 NAND2X1_1285 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n149), .Y(reg_ve__abc_3798_n150) );
	NAND2X1 NAND2X1_1286 ( .A(reset), .B(vdd), .Y(reg_ve__abc_3798_n151) );
	NAND2X1 NAND2X1_1287 ( .A(reg_ve__abc_3798_n151), .B(reg_ve__abc_3798_n150), .Y(reg_ve_value_2__FF_INPUT) );
	NOR2X1 NOR2X1_815 ( .A(reset), .B(reg_ve__abc_3798_n96), .Y(reg_ve__abc_3798_n153) );
	NAND2X1 NAND2X1_1288 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n153), .Y(reg_ve__abc_3798_n154) );
	NAND2X1 NAND2X1_1289 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n155) );
	NAND2X1 NAND2X1_1290 ( .A(reg_ve__abc_3798_n155), .B(reg_ve__abc_3798_n154), .Y(reg_ve__abc_3798_n74) );
	NOR2X1 NOR2X1_816 ( .A(reset), .B(reg_ve__abc_3798_n98), .Y(reg_ve__abc_3798_n157) );
	NAND2X1 NAND2X1_1291 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n157), .Y(reg_ve__abc_3798_n158) );
	NAND2X1 NAND2X1_1292 ( .A(reset), .B(vdd), .Y(reg_ve__abc_3798_n159) );
	NAND2X1 NAND2X1_1293 ( .A(reg_ve__abc_3798_n159), .B(reg_ve__abc_3798_n158), .Y(reg_ve_value_0__FF_INPUT) );
	INVX1 INVX1_339 ( .A(reg_ve_value_15_), .Y(reg_ve__abc_3798_n161) );
	NOR2X1 NOR2X1_817 ( .A(reset), .B(reg_ve__abc_3798_n161), .Y(reg_ve__abc_3798_n162) );
	NAND2X1 NAND2X1_1294 ( .A(reg_ve__abc_3798_n100), .B(reg_ve__abc_3798_n162), .Y(reg_ve__abc_3798_n163) );
	NAND2X1 NAND2X1_1295 ( .A(reset), .B(gnd), .Y(reg_ve__abc_3798_n164) );
	NAND2X1 NAND2X1_1296 ( .A(reg_ve__abc_3798_n164), .B(reg_ve__abc_3798_n163), .Y(reg_ve_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_818 ( .A(reg_ve__abc_3798_n161), .B(reg_ve__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_258 ( .CLK(clk), .D(reg_ve_value_0__FF_INPUT), .Q(reg_ve_value_0_) );
	DFFPOSX1 DFFPOSX1_259 ( .CLK(clk), .D(reg_ve__abc_3798_n74), .Q(reg_ve_value_1_) );
	DFFPOSX1 DFFPOSX1_260 ( .CLK(clk), .D(reg_ve_value_2__FF_INPUT), .Q(reg_ve_value_2_) );
	DFFPOSX1 DFFPOSX1_261 ( .CLK(clk), .D(reg_ve_value_3__FF_INPUT), .Q(reg_ve_value_3_) );
	DFFPOSX1 DFFPOSX1_262 ( .CLK(clk), .D(reg_ve__abc_3798_n65), .Q(reg_ve_value_4_) );
	DFFPOSX1 DFFPOSX1_263 ( .CLK(clk), .D(reg_ve_value_5__FF_INPUT), .Q(reg_ve_value_5_) );
	DFFPOSX1 DFFPOSX1_264 ( .CLK(clk), .D(reg_ve_value_6__FF_INPUT), .Q(reg_ve_value_6_) );
	DFFPOSX1 DFFPOSX1_265 ( .CLK(clk), .D(reg_ve__abc_3798_n56), .Q(reg_ve_value_7_) );
	DFFPOSX1 DFFPOSX1_266 ( .CLK(clk), .D(reg_ve__abc_3798_n53), .Q(reg_ve_value_8_) );
	DFFPOSX1 DFFPOSX1_267 ( .CLK(clk), .D(reg_ve_value_9__FF_INPUT), .Q(reg_ve_value_9_) );
	DFFPOSX1 DFFPOSX1_268 ( .CLK(clk), .D(reg_ve__abc_3798_n47), .Q(reg_ve_value_10_) );
	DFFPOSX1 DFFPOSX1_269 ( .CLK(clk), .D(reg_ve__abc_3798_n44), .Q(reg_ve_value_11_) );
	DFFPOSX1 DFFPOSX1_270 ( .CLK(clk), .D(reg_ve_value_12__FF_INPUT), .Q(reg_ve_value_12_) );
	DFFPOSX1 DFFPOSX1_271 ( .CLK(clk), .D(reg_ve_value_13__FF_INPUT), .Q(reg_ve_value_13_) );
	DFFPOSX1 DFFPOSX1_272 ( .CLK(clk), .D(reg_ve__abc_3798_n35), .Q(reg_ve_value_14_) );
	DFFPOSX1 DFFPOSX1_273 ( .CLK(clk), .D(reg_ve_value_15__FF_INPUT), .Q(reg_ve_value_15_) );
	INVX1 INVX1_340 ( .A(reg_vf_value_14_), .Y(reg_vf__abc_3798_n68_1) );
	INVX1 INVX1_341 ( .A(we), .Y(reg_vf__abc_3798_n69) );
	NAND2X1 NAND2X1_1297 ( .A(addr_vf), .B(reg_vf__abc_3798_n69), .Y(reg_vf__abc_3798_n70_1) );
	NOR2X1 NOR2X1_819 ( .A(reg_vf__abc_3798_n68_1), .B(reg_vf__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_342 ( .A(reg_vf_value_13_), .Y(reg_vf__abc_3798_n72) );
	NOR2X1 NOR2X1_820 ( .A(reg_vf__abc_3798_n72), .B(reg_vf__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_343 ( .A(reg_vf_value_12_), .Y(reg_vf__abc_3798_n74_1) );
	NOR2X1 NOR2X1_821 ( .A(reg_vf__abc_3798_n74_1), .B(reg_vf__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_344 ( .A(reg_vf_value_11_), .Y(reg_vf__abc_3798_n76_1) );
	NOR2X1 NOR2X1_822 ( .A(reg_vf__abc_3798_n76_1), .B(reg_vf__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_345 ( .A(reg_vf_value_10_), .Y(reg_vf__abc_3798_n78) );
	NOR2X1 NOR2X1_823 ( .A(reg_vf__abc_3798_n78), .B(reg_vf__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_346 ( .A(reg_vf_value_9_), .Y(reg_vf__abc_3798_n80_1) );
	NOR2X1 NOR2X1_824 ( .A(reg_vf__abc_3798_n80_1), .B(reg_vf__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_347 ( .A(reg_vf_value_8_), .Y(reg_vf__abc_3798_n82_1) );
	NOR2X1 NOR2X1_825 ( .A(reg_vf__abc_3798_n82_1), .B(reg_vf__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_348 ( .A(reg_vf_value_7_), .Y(reg_vf__abc_3798_n84_1) );
	NOR2X1 NOR2X1_826 ( .A(reg_vf__abc_3798_n84_1), .B(reg_vf__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_349 ( .A(reg_vf_value_6_), .Y(reg_vf__abc_3798_n86) );
	NOR2X1 NOR2X1_827 ( .A(reg_vf__abc_3798_n86), .B(reg_vf__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_350 ( .A(reg_vf_value_5_), .Y(reg_vf__abc_3798_n88) );
	NOR2X1 NOR2X1_828 ( .A(reg_vf__abc_3798_n88), .B(reg_vf__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_351 ( .A(reg_vf_value_4_), .Y(reg_vf__abc_3798_n90) );
	NOR2X1 NOR2X1_829 ( .A(reg_vf__abc_3798_n90), .B(reg_vf__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_352 ( .A(reg_vf_value_3_), .Y(reg_vf__abc_3798_n92) );
	NOR2X1 NOR2X1_830 ( .A(reg_vf__abc_3798_n92), .B(reg_vf__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_353 ( .A(reg_vf_value_2_), .Y(reg_vf__abc_3798_n94) );
	NOR2X1 NOR2X1_831 ( .A(reg_vf__abc_3798_n94), .B(reg_vf__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_354 ( .A(reg_vf_value_1_), .Y(reg_vf__abc_3798_n96) );
	NOR2X1 NOR2X1_832 ( .A(reg_vf__abc_3798_n96), .B(reg_vf__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_355 ( .A(reg_vf_value_0_), .Y(reg_vf__abc_3798_n98) );
	NOR2X1 NOR2X1_833 ( .A(reg_vf__abc_3798_n98), .B(reg_vf__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1298 ( .A(we), .B(addr_vf), .Y(reg_vf__abc_3798_n100) );
	NOR2X1 NOR2X1_834 ( .A(reset), .B(reg_vf__abc_3798_n68_1), .Y(reg_vf__abc_3798_n101) );
	NAND2X1 NAND2X1_1299 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n101), .Y(reg_vf__abc_3798_n102) );
	NAND2X1 NAND2X1_1300 ( .A(gnd), .B(reset), .Y(reg_vf__abc_3798_n103) );
	NAND2X1 NAND2X1_1301 ( .A(reg_vf__abc_3798_n103), .B(reg_vf__abc_3798_n102), .Y(reg_vf_value_14__FF_INPUT) );
	NOR2X1 NOR2X1_835 ( .A(reset), .B(reg_vf__abc_3798_n72), .Y(reg_vf__abc_3798_n105) );
	NAND2X1 NAND2X1_1302 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n105), .Y(reg_vf__abc_3798_n106) );
	NAND2X1 NAND2X1_1303 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n107) );
	NAND2X1 NAND2X1_1304 ( .A(reg_vf__abc_3798_n107), .B(reg_vf__abc_3798_n106), .Y(reg_vf__abc_3798_n38) );
	NOR2X1 NOR2X1_836 ( .A(reset), .B(reg_vf__abc_3798_n74_1), .Y(reg_vf__abc_3798_n109) );
	NAND2X1 NAND2X1_1305 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n109), .Y(reg_vf__abc_3798_n110) );
	NAND2X1 NAND2X1_1306 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n111) );
	NAND2X1 NAND2X1_1307 ( .A(reg_vf__abc_3798_n111), .B(reg_vf__abc_3798_n110), .Y(reg_vf_value_12__FF_INPUT) );
	NOR2X1 NOR2X1_837 ( .A(reset), .B(reg_vf__abc_3798_n76_1), .Y(reg_vf__abc_3798_n113) );
	NAND2X1 NAND2X1_1308 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n113), .Y(reg_vf__abc_3798_n114) );
	NAND2X1 NAND2X1_1309 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n115) );
	NAND2X1 NAND2X1_1310 ( .A(reg_vf__abc_3798_n115), .B(reg_vf__abc_3798_n114), .Y(reg_vf__abc_3798_n44) );
	NOR2X1 NOR2X1_838 ( .A(reset), .B(reg_vf__abc_3798_n78), .Y(reg_vf__abc_3798_n117) );
	NAND2X1 NAND2X1_1311 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n117), .Y(reg_vf__abc_3798_n118) );
	NAND2X1 NAND2X1_1312 ( .A(reset), .B(vdd), .Y(reg_vf__abc_3798_n119) );
	NAND2X1 NAND2X1_1313 ( .A(reg_vf__abc_3798_n119), .B(reg_vf__abc_3798_n118), .Y(reg_vf__abc_3798_n47) );
	NOR2X1 NOR2X1_839 ( .A(reset), .B(reg_vf__abc_3798_n80_1), .Y(reg_vf__abc_3798_n121) );
	NAND2X1 NAND2X1_1314 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n121), .Y(reg_vf__abc_3798_n122) );
	NAND2X1 NAND2X1_1315 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n123) );
	NAND2X1 NAND2X1_1316 ( .A(reg_vf__abc_3798_n123), .B(reg_vf__abc_3798_n122), .Y(reg_vf_value_9__FF_INPUT) );
	NOR2X1 NOR2X1_840 ( .A(reset), .B(reg_vf__abc_3798_n82_1), .Y(reg_vf__abc_3798_n125) );
	NAND2X1 NAND2X1_1317 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n125), .Y(reg_vf__abc_3798_n126) );
	NAND2X1 NAND2X1_1318 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n127) );
	NAND2X1 NAND2X1_1319 ( .A(reg_vf__abc_3798_n127), .B(reg_vf__abc_3798_n126), .Y(reg_vf_value_8__FF_INPUT) );
	NOR2X1 NOR2X1_841 ( .A(reset), .B(reg_vf__abc_3798_n84_1), .Y(reg_vf__abc_3798_n129) );
	NAND2X1 NAND2X1_1320 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n129), .Y(reg_vf__abc_3798_n130) );
	NAND2X1 NAND2X1_1321 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n131) );
	NAND2X1 NAND2X1_1322 ( .A(reg_vf__abc_3798_n131), .B(reg_vf__abc_3798_n130), .Y(reg_vf__abc_3798_n56) );
	NOR2X1 NOR2X1_842 ( .A(reset), .B(reg_vf__abc_3798_n86), .Y(reg_vf__abc_3798_n133) );
	NAND2X1 NAND2X1_1323 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n133), .Y(reg_vf__abc_3798_n134) );
	NAND2X1 NAND2X1_1324 ( .A(reset), .B(vdd), .Y(reg_vf__abc_3798_n135) );
	NAND2X1 NAND2X1_1325 ( .A(reg_vf__abc_3798_n135), .B(reg_vf__abc_3798_n134), .Y(reg_vf_value_6__FF_INPUT) );
	NOR2X1 NOR2X1_843 ( .A(reset), .B(reg_vf__abc_3798_n88), .Y(reg_vf__abc_3798_n137) );
	NAND2X1 NAND2X1_1326 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n137), .Y(reg_vf__abc_3798_n138) );
	NAND2X1 NAND2X1_1327 ( .A(reset), .B(vdd), .Y(reg_vf__abc_3798_n139) );
	NAND2X1 NAND2X1_1328 ( .A(reg_vf__abc_3798_n139), .B(reg_vf__abc_3798_n138), .Y(reg_vf__abc_3798_n62) );
	NOR2X1 NOR2X1_844 ( .A(reset), .B(reg_vf__abc_3798_n90), .Y(reg_vf__abc_3798_n141) );
	NAND2X1 NAND2X1_1329 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n141), .Y(reg_vf__abc_3798_n142) );
	NAND2X1 NAND2X1_1330 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n143) );
	NAND2X1 NAND2X1_1331 ( .A(reg_vf__abc_3798_n143), .B(reg_vf__abc_3798_n142), .Y(reg_vf__abc_3798_n65) );
	NOR2X1 NOR2X1_845 ( .A(reset), .B(reg_vf__abc_3798_n92), .Y(reg_vf__abc_3798_n145) );
	NAND2X1 NAND2X1_1332 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n145), .Y(reg_vf__abc_3798_n146) );
	NAND2X1 NAND2X1_1333 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n147) );
	NAND2X1 NAND2X1_1334 ( .A(reg_vf__abc_3798_n147), .B(reg_vf__abc_3798_n146), .Y(reg_vf_value_3__FF_INPUT) );
	NOR2X1 NOR2X1_846 ( .A(reset), .B(reg_vf__abc_3798_n94), .Y(reg_vf__abc_3798_n149) );
	NAND2X1 NAND2X1_1335 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n149), .Y(reg_vf__abc_3798_n150) );
	NAND2X1 NAND2X1_1336 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n151) );
	NAND2X1 NAND2X1_1337 ( .A(reg_vf__abc_3798_n151), .B(reg_vf__abc_3798_n150), .Y(reg_vf__abc_3798_n71) );
	NOR2X1 NOR2X1_847 ( .A(reset), .B(reg_vf__abc_3798_n96), .Y(reg_vf__abc_3798_n153) );
	NAND2X1 NAND2X1_1338 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n153), .Y(reg_vf__abc_3798_n154) );
	NAND2X1 NAND2X1_1339 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n155) );
	NAND2X1 NAND2X1_1340 ( .A(reg_vf__abc_3798_n155), .B(reg_vf__abc_3798_n154), .Y(reg_vf__abc_3798_n74) );
	NOR2X1 NOR2X1_848 ( .A(reset), .B(reg_vf__abc_3798_n98), .Y(reg_vf__abc_3798_n157) );
	NAND2X1 NAND2X1_1341 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n157), .Y(reg_vf__abc_3798_n158) );
	NAND2X1 NAND2X1_1342 ( .A(reset), .B(vdd), .Y(reg_vf__abc_3798_n159) );
	NAND2X1 NAND2X1_1343 ( .A(reg_vf__abc_3798_n159), .B(reg_vf__abc_3798_n158), .Y(reg_vf__abc_3798_n77) );
	INVX1 INVX1_356 ( .A(reg_vf_value_15_), .Y(reg_vf__abc_3798_n161) );
	NOR2X1 NOR2X1_849 ( .A(reset), .B(reg_vf__abc_3798_n161), .Y(reg_vf__abc_3798_n162) );
	NAND2X1 NAND2X1_1344 ( .A(reg_vf__abc_3798_n100), .B(reg_vf__abc_3798_n162), .Y(reg_vf__abc_3798_n163) );
	NAND2X1 NAND2X1_1345 ( .A(reset), .B(gnd), .Y(reg_vf__abc_3798_n164) );
	NAND2X1 NAND2X1_1346 ( .A(reg_vf__abc_3798_n164), .B(reg_vf__abc_3798_n163), .Y(reg_vf_value_15__FF_INPUT) );
	NOR2X1 NOR2X1_850 ( .A(reg_vf__abc_3798_n161), .B(reg_vf__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_274 ( .CLK(clk), .D(reg_vf__abc_3798_n77), .Q(reg_vf_value_0_) );
	DFFPOSX1 DFFPOSX1_275 ( .CLK(clk), .D(reg_vf__abc_3798_n74), .Q(reg_vf_value_1_) );
	DFFPOSX1 DFFPOSX1_276 ( .CLK(clk), .D(reg_vf__abc_3798_n71), .Q(reg_vf_value_2_) );
	DFFPOSX1 DFFPOSX1_277 ( .CLK(clk), .D(reg_vf_value_3__FF_INPUT), .Q(reg_vf_value_3_) );
	DFFPOSX1 DFFPOSX1_278 ( .CLK(clk), .D(reg_vf__abc_3798_n65), .Q(reg_vf_value_4_) );
	DFFPOSX1 DFFPOSX1_279 ( .CLK(clk), .D(reg_vf__abc_3798_n62), .Q(reg_vf_value_5_) );
	DFFPOSX1 DFFPOSX1_280 ( .CLK(clk), .D(reg_vf_value_6__FF_INPUT), .Q(reg_vf_value_6_) );
	DFFPOSX1 DFFPOSX1_281 ( .CLK(clk), .D(reg_vf__abc_3798_n56), .Q(reg_vf_value_7_) );
	DFFPOSX1 DFFPOSX1_282 ( .CLK(clk), .D(reg_vf_value_8__FF_INPUT), .Q(reg_vf_value_8_) );
	DFFPOSX1 DFFPOSX1_283 ( .CLK(clk), .D(reg_vf_value_9__FF_INPUT), .Q(reg_vf_value_9_) );
	DFFPOSX1 DFFPOSX1_284 ( .CLK(clk), .D(reg_vf__abc_3798_n47), .Q(reg_vf_value_10_) );
	DFFPOSX1 DFFPOSX1_285 ( .CLK(clk), .D(reg_vf__abc_3798_n44), .Q(reg_vf_value_11_) );
	DFFPOSX1 DFFPOSX1_286 ( .CLK(clk), .D(reg_vf_value_12__FF_INPUT), .Q(reg_vf_value_12_) );
	DFFPOSX1 DFFPOSX1_287 ( .CLK(clk), .D(reg_vf__abc_3798_n38), .Q(reg_vf_value_13_) );
	DFFPOSX1 DFFPOSX1_288 ( .CLK(clk), .D(reg_vf_value_14__FF_INPUT), .Q(reg_vf_value_14_) );
	DFFPOSX1 DFFPOSX1_289 ( .CLK(clk), .D(reg_vf_value_15__FF_INPUT), .Q(reg_vf_value_15_) );
	INVX1 INVX1_357 ( .A(reg_vv_value_14_), .Y(reg_vv__abc_3798_n68_1) );
	INVX1 INVX1_358 ( .A(we), .Y(reg_vv__abc_3798_n69) );
	NAND2X1 NAND2X1_1347 ( .A(addr_vv), .B(reg_vv__abc_3798_n69), .Y(reg_vv__abc_3798_n70_1) );
	NOR2X1 NOR2X1_851 ( .A(reg_vv__abc_3798_n68_1), .B(reg_vv__abc_3798_n70_1), .Y(data[14]) );
	INVX1 INVX1_359 ( .A(reg_vv_value_13_), .Y(reg_vv__abc_3798_n72) );
	NOR2X1 NOR2X1_852 ( .A(reg_vv__abc_3798_n72), .B(reg_vv__abc_3798_n70_1), .Y(data[13]) );
	INVX1 INVX1_360 ( .A(reg_vv_value_12_), .Y(reg_vv__abc_3798_n74_1) );
	NOR2X1 NOR2X1_853 ( .A(reg_vv__abc_3798_n74_1), .B(reg_vv__abc_3798_n70_1), .Y(data[12]) );
	INVX1 INVX1_361 ( .A(reg_vv_value_11_), .Y(reg_vv__abc_3798_n76_1) );
	NOR2X1 NOR2X1_854 ( .A(reg_vv__abc_3798_n76_1), .B(reg_vv__abc_3798_n70_1), .Y(data[11]) );
	INVX1 INVX1_362 ( .A(reg_vv_value_10_), .Y(reg_vv__abc_3798_n78) );
	NOR2X1 NOR2X1_855 ( .A(reg_vv__abc_3798_n78), .B(reg_vv__abc_3798_n70_1), .Y(data[10]) );
	INVX1 INVX1_363 ( .A(reg_vv_value_9_), .Y(reg_vv__abc_3798_n80_1) );
	NOR2X1 NOR2X1_856 ( .A(reg_vv__abc_3798_n80_1), .B(reg_vv__abc_3798_n70_1), .Y(data[9]) );
	INVX1 INVX1_364 ( .A(reg_vv_value_8_), .Y(reg_vv__abc_3798_n82_1) );
	NOR2X1 NOR2X1_857 ( .A(reg_vv__abc_3798_n82_1), .B(reg_vv__abc_3798_n70_1), .Y(data[8]) );
	INVX1 INVX1_365 ( .A(reg_vv_value_7_), .Y(reg_vv__abc_3798_n84_1) );
	NOR2X1 NOR2X1_858 ( .A(reg_vv__abc_3798_n84_1), .B(reg_vv__abc_3798_n70_1), .Y(data[7]) );
	INVX1 INVX1_366 ( .A(reg_vv_value_6_), .Y(reg_vv__abc_3798_n86) );
	NOR2X1 NOR2X1_859 ( .A(reg_vv__abc_3798_n86), .B(reg_vv__abc_3798_n70_1), .Y(data[6]) );
	INVX1 INVX1_367 ( .A(reg_vv_value_5_), .Y(reg_vv__abc_3798_n88) );
	NOR2X1 NOR2X1_860 ( .A(reg_vv__abc_3798_n88), .B(reg_vv__abc_3798_n70_1), .Y(data[5]) );
	INVX1 INVX1_368 ( .A(reg_vv_value_4_), .Y(reg_vv__abc_3798_n90) );
	NOR2X1 NOR2X1_861 ( .A(reg_vv__abc_3798_n90), .B(reg_vv__abc_3798_n70_1), .Y(data[4]) );
	INVX1 INVX1_369 ( .A(reg_vv_value_3_), .Y(reg_vv__abc_3798_n92) );
	NOR2X1 NOR2X1_862 ( .A(reg_vv__abc_3798_n92), .B(reg_vv__abc_3798_n70_1), .Y(data[3]) );
	INVX1 INVX1_370 ( .A(reg_vv_value_2_), .Y(reg_vv__abc_3798_n94) );
	NOR2X1 NOR2X1_863 ( .A(reg_vv__abc_3798_n94), .B(reg_vv__abc_3798_n70_1), .Y(data[2]) );
	INVX1 INVX1_371 ( .A(reg_vv_value_1_), .Y(reg_vv__abc_3798_n96) );
	NOR2X1 NOR2X1_864 ( .A(reg_vv__abc_3798_n96), .B(reg_vv__abc_3798_n70_1), .Y(data[1]) );
	INVX1 INVX1_372 ( .A(reg_vv_value_0_), .Y(reg_vv__abc_3798_n98) );
	NOR2X1 NOR2X1_865 ( .A(reg_vv__abc_3798_n98), .B(reg_vv__abc_3798_n70_1), .Y(data[0]) );
	NAND2X1 NAND2X1_1348 ( .A(we), .B(addr_vv), .Y(reg_vv__abc_3798_n100) );
	NOR2X1 NOR2X1_866 ( .A(reset), .B(reg_vv__abc_3798_n68_1), .Y(reg_vv__abc_3798_n101) );
	NAND2X1 NAND2X1_1349 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n101), .Y(reg_vv__abc_3798_n102) );
	NAND2X1 NAND2X1_1350 ( .A(gnd), .B(reset), .Y(reg_vv__abc_3798_n103) );
	NAND2X1 NAND2X1_1351 ( .A(reg_vv__abc_3798_n103), .B(reg_vv__abc_3798_n102), .Y(reg_vv__abc_3798_n35) );
	NOR2X1 NOR2X1_867 ( .A(reset), .B(reg_vv__abc_3798_n72), .Y(reg_vv__abc_3798_n105) );
	NAND2X1 NAND2X1_1352 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n105), .Y(reg_vv__abc_3798_n106) );
	NAND2X1 NAND2X1_1353 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n107) );
	NAND2X1 NAND2X1_1354 ( .A(reg_vv__abc_3798_n107), .B(reg_vv__abc_3798_n106), .Y(reg_vv__abc_3798_n38) );
	NOR2X1 NOR2X1_868 ( .A(reset), .B(reg_vv__abc_3798_n74_1), .Y(reg_vv__abc_3798_n109) );
	NAND2X1 NAND2X1_1355 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n109), .Y(reg_vv__abc_3798_n110) );
	NAND2X1 NAND2X1_1356 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n111) );
	NAND2X1 NAND2X1_1357 ( .A(reg_vv__abc_3798_n111), .B(reg_vv__abc_3798_n110), .Y(reg_vv__abc_3798_n41) );
	NOR2X1 NOR2X1_869 ( .A(reset), .B(reg_vv__abc_3798_n76_1), .Y(reg_vv__abc_3798_n113) );
	NAND2X1 NAND2X1_1358 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n113), .Y(reg_vv__abc_3798_n114) );
	NAND2X1 NAND2X1_1359 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n115) );
	NAND2X1 NAND2X1_1360 ( .A(reg_vv__abc_3798_n115), .B(reg_vv__abc_3798_n114), .Y(reg_vv__abc_3798_n44) );
	NOR2X1 NOR2X1_870 ( .A(reset), .B(reg_vv__abc_3798_n78), .Y(reg_vv__abc_3798_n117) );
	NAND2X1 NAND2X1_1361 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n117), .Y(reg_vv__abc_3798_n118) );
	NAND2X1 NAND2X1_1362 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n119) );
	NAND2X1 NAND2X1_1363 ( .A(reg_vv__abc_3798_n119), .B(reg_vv__abc_3798_n118), .Y(reg_vv__abc_3798_n47) );
	NOR2X1 NOR2X1_871 ( .A(reset), .B(reg_vv__abc_3798_n80_1), .Y(reg_vv__abc_3798_n121) );
	NAND2X1 NAND2X1_1364 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n121), .Y(reg_vv__abc_3798_n122) );
	NAND2X1 NAND2X1_1365 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n123) );
	NAND2X1 NAND2X1_1366 ( .A(reg_vv__abc_3798_n123), .B(reg_vv__abc_3798_n122), .Y(reg_vv__abc_3798_n50) );
	NOR2X1 NOR2X1_872 ( .A(reset), .B(reg_vv__abc_3798_n82_1), .Y(reg_vv__abc_3798_n125) );
	NAND2X1 NAND2X1_1367 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n125), .Y(reg_vv__abc_3798_n126) );
	NAND2X1 NAND2X1_1368 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n127) );
	NAND2X1 NAND2X1_1369 ( .A(reg_vv__abc_3798_n127), .B(reg_vv__abc_3798_n126), .Y(reg_vv__abc_3798_n53) );
	NOR2X1 NOR2X1_873 ( .A(reset), .B(reg_vv__abc_3798_n84_1), .Y(reg_vv__abc_3798_n129) );
	NAND2X1 NAND2X1_1370 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n129), .Y(reg_vv__abc_3798_n130) );
	NAND2X1 NAND2X1_1371 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n131) );
	NAND2X1 NAND2X1_1372 ( .A(reg_vv__abc_3798_n131), .B(reg_vv__abc_3798_n130), .Y(reg_vv__abc_3798_n56) );
	NOR2X1 NOR2X1_874 ( .A(reset), .B(reg_vv__abc_3798_n86), .Y(reg_vv__abc_3798_n133) );
	NAND2X1 NAND2X1_1373 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n133), .Y(reg_vv__abc_3798_n134) );
	NAND2X1 NAND2X1_1374 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n135) );
	NAND2X1 NAND2X1_1375 ( .A(reg_vv__abc_3798_n135), .B(reg_vv__abc_3798_n134), .Y(reg_vv__abc_3798_n59) );
	NOR2X1 NOR2X1_875 ( .A(reset), .B(reg_vv__abc_3798_n88), .Y(reg_vv__abc_3798_n137) );
	NAND2X1 NAND2X1_1376 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n137), .Y(reg_vv__abc_3798_n138) );
	NAND2X1 NAND2X1_1377 ( .A(reset), .B(vdd), .Y(reg_vv__abc_3798_n139) );
	NAND2X1 NAND2X1_1378 ( .A(reg_vv__abc_3798_n139), .B(reg_vv__abc_3798_n138), .Y(reg_vv__abc_3798_n62) );
	NOR2X1 NOR2X1_876 ( .A(reset), .B(reg_vv__abc_3798_n90), .Y(reg_vv__abc_3798_n141) );
	NAND2X1 NAND2X1_1379 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n141), .Y(reg_vv__abc_3798_n142) );
	NAND2X1 NAND2X1_1380 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n143) );
	NAND2X1 NAND2X1_1381 ( .A(reg_vv__abc_3798_n143), .B(reg_vv__abc_3798_n142), .Y(reg_vv__abc_3798_n65) );
	NOR2X1 NOR2X1_877 ( .A(reset), .B(reg_vv__abc_3798_n92), .Y(reg_vv__abc_3798_n145) );
	NAND2X1 NAND2X1_1382 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n145), .Y(reg_vv__abc_3798_n146) );
	NAND2X1 NAND2X1_1383 ( .A(reset), .B(vdd), .Y(reg_vv__abc_3798_n147) );
	NAND2X1 NAND2X1_1384 ( .A(reg_vv__abc_3798_n147), .B(reg_vv__abc_3798_n146), .Y(reg_vv__abc_3798_n68) );
	NOR2X1 NOR2X1_878 ( .A(reset), .B(reg_vv__abc_3798_n94), .Y(reg_vv__abc_3798_n149) );
	NAND2X1 NAND2X1_1385 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n149), .Y(reg_vv__abc_3798_n150) );
	NAND2X1 NAND2X1_1386 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n151) );
	NAND2X1 NAND2X1_1387 ( .A(reg_vv__abc_3798_n151), .B(reg_vv__abc_3798_n150), .Y(reg_vv__abc_3798_n71) );
	NOR2X1 NOR2X1_879 ( .A(reset), .B(reg_vv__abc_3798_n96), .Y(reg_vv__abc_3798_n153) );
	NAND2X1 NAND2X1_1388 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n153), .Y(reg_vv__abc_3798_n154) );
	NAND2X1 NAND2X1_1389 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n155) );
	NAND2X1 NAND2X1_1390 ( .A(reg_vv__abc_3798_n155), .B(reg_vv__abc_3798_n154), .Y(reg_vv__abc_3798_n74) );
	NOR2X1 NOR2X1_880 ( .A(reset), .B(reg_vv__abc_3798_n98), .Y(reg_vv__abc_3798_n157) );
	NAND2X1 NAND2X1_1391 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n157), .Y(reg_vv__abc_3798_n158) );
	NAND2X1 NAND2X1_1392 ( .A(reset), .B(vdd), .Y(reg_vv__abc_3798_n159) );
	NAND2X1 NAND2X1_1393 ( .A(reg_vv__abc_3798_n159), .B(reg_vv__abc_3798_n158), .Y(reg_vv__abc_3798_n77) );
	INVX1 INVX1_373 ( .A(reg_vv_value_15_), .Y(reg_vv__abc_3798_n161) );
	NOR2X1 NOR2X1_881 ( .A(reset), .B(reg_vv__abc_3798_n161), .Y(reg_vv__abc_3798_n162) );
	NAND2X1 NAND2X1_1394 ( .A(reg_vv__abc_3798_n100), .B(reg_vv__abc_3798_n162), .Y(reg_vv__abc_3798_n163) );
	NAND2X1 NAND2X1_1395 ( .A(reset), .B(gnd), .Y(reg_vv__abc_3798_n164) );
	NAND2X1 NAND2X1_1396 ( .A(reg_vv__abc_3798_n164), .B(reg_vv__abc_3798_n163), .Y(reg_vv__abc_3798_n81) );
	NOR2X1 NOR2X1_882 ( .A(reg_vv__abc_3798_n161), .B(reg_vv__abc_3798_n70_1), .Y(data[15]) );
	DFFPOSX1 DFFPOSX1_290 ( .CLK(clk), .D(reg_vv__abc_3798_n77), .Q(reg_vv_value_0_) );
	DFFPOSX1 DFFPOSX1_291 ( .CLK(clk), .D(reg_vv__abc_3798_n74), .Q(reg_vv_value_1_) );
	DFFPOSX1 DFFPOSX1_292 ( .CLK(clk), .D(reg_vv__abc_3798_n71), .Q(reg_vv_value_2_) );
	DFFPOSX1 DFFPOSX1_293 ( .CLK(clk), .D(reg_vv__abc_3798_n68), .Q(reg_vv_value_3_) );
	DFFPOSX1 DFFPOSX1_294 ( .CLK(clk), .D(reg_vv__abc_3798_n65), .Q(reg_vv_value_4_) );
	DFFPOSX1 DFFPOSX1_295 ( .CLK(clk), .D(reg_vv__abc_3798_n62), .Q(reg_vv_value_5_) );
	DFFPOSX1 DFFPOSX1_296 ( .CLK(clk), .D(reg_vv__abc_3798_n59), .Q(reg_vv_value_6_) );
	DFFPOSX1 DFFPOSX1_297 ( .CLK(clk), .D(reg_vv__abc_3798_n56), .Q(reg_vv_value_7_) );
	DFFPOSX1 DFFPOSX1_298 ( .CLK(clk), .D(reg_vv__abc_3798_n53), .Q(reg_vv_value_8_) );
	DFFPOSX1 DFFPOSX1_299 ( .CLK(clk), .D(reg_vv__abc_3798_n50), .Q(reg_vv_value_9_) );
	DFFPOSX1 DFFPOSX1_300 ( .CLK(clk), .D(reg_vv__abc_3798_n47), .Q(reg_vv_value_10_) );
	DFFPOSX1 DFFPOSX1_301 ( .CLK(clk), .D(reg_vv__abc_3798_n44), .Q(reg_vv_value_11_) );
	DFFPOSX1 DFFPOSX1_302 ( .CLK(clk), .D(reg_vv__abc_3798_n41), .Q(reg_vv_value_12_) );
	DFFPOSX1 DFFPOSX1_303 ( .CLK(clk), .D(reg_vv__abc_3798_n38), .Q(reg_vv_value_13_) );
	DFFPOSX1 DFFPOSX1_304 ( .CLK(clk), .D(reg_vv__abc_3798_n35), .Q(reg_vv_value_14_) );
	DFFPOSX1 DFFPOSX1_305 ( .CLK(clk), .D(reg_vv__abc_3798_n81), .Q(reg_vv_value_15_) );
	BUFX2 BUFX2_40 ( .A(clk), .Y(reg_sh_clk) );
	BUFX2 BUFX2_41 ( .A(reset), .Y(reg_sh_reset) );
	BUFX2 BUFX2_42 ( .A(addr_sh), .Y(reg_sh_cs) );
	BUFX2 BUFX2_43 ( .A(we), .Y(reg_sh_we) );
	BUFX2 BUFX2_44 ( .A(data[0]), .Y(reg_sh_data_0_) );
	BUFX2 BUFX2_45 ( .A(data[1]), .Y(reg_sh_data_1_) );
	BUFX2 BUFX2_46 ( .A(data[2]), .Y(reg_sh_data_2_) );
	BUFX2 BUFX2_47 ( .A(data[3]), .Y(reg_sh_data_3_) );
	BUFX2 BUFX2_48 ( .A(data[4]), .Y(reg_sh_data_4_) );
	BUFX2 BUFX2_49 ( .A(data[5]), .Y(reg_sh_data_5_) );
	BUFX2 BUFX2_50 ( .A(data[6]), .Y(reg_sh_data_6_) );
	BUFX2 BUFX2_51 ( .A(data[7]), .Y(reg_sh_data_7_) );
	BUFX2 BUFX2_52 ( .A(data[8]), .Y(reg_sh_data_8_) );
	BUFX2 BUFX2_53 ( .A(data[9]), .Y(reg_sh_data_9_) );
	BUFX2 BUFX2_54 ( .A(data[10]), .Y(reg_sh_data_10_) );
	BUFX2 BUFX2_55 ( .A(data[11]), .Y(reg_sh_data_11_) );
	BUFX2 BUFX2_56 ( .A(data[12]), .Y(reg_sh_data_12_) );
	BUFX2 BUFX2_57 ( .A(data[13]), .Y(reg_sh_data_13_) );
	BUFX2 BUFX2_58 ( .A(data[14]), .Y(reg_sh_data_14_) );
	BUFX2 BUFX2_59 ( .A(data[15]), .Y(reg_sh_data_15_) );
	BUFX2 BUFX2_60 ( .A(clk), .Y(reg_fl_clk) );
	BUFX2 BUFX2_61 ( .A(reset), .Y(reg_fl_reset) );
	BUFX2 BUFX2_62 ( .A(addr_fl), .Y(reg_fl_cs) );
	BUFX2 BUFX2_63 ( .A(we), .Y(reg_fl_we) );
	BUFX2 BUFX2_64 ( .A(data[0]), .Y(reg_fl_data_0_) );
	BUFX2 BUFX2_65 ( .A(data[1]), .Y(reg_fl_data_1_) );
	BUFX2 BUFX2_66 ( .A(data[2]), .Y(reg_fl_data_2_) );
	BUFX2 BUFX2_67 ( .A(data[3]), .Y(reg_fl_data_3_) );
	BUFX2 BUFX2_68 ( .A(data[4]), .Y(reg_fl_data_4_) );
	BUFX2 BUFX2_69 ( .A(data[5]), .Y(reg_fl_data_5_) );
	BUFX2 BUFX2_70 ( .A(data[6]), .Y(reg_fl_data_6_) );
	BUFX2 BUFX2_71 ( .A(data[7]), .Y(reg_fl_data_7_) );
	BUFX2 BUFX2_72 ( .A(data[8]), .Y(reg_fl_data_8_) );
	BUFX2 BUFX2_73 ( .A(data[9]), .Y(reg_fl_data_9_) );
	BUFX2 BUFX2_74 ( .A(data[10]), .Y(reg_fl_data_10_) );
	BUFX2 BUFX2_75 ( .A(data[11]), .Y(reg_fl_data_11_) );
	BUFX2 BUFX2_76 ( .A(data[12]), .Y(reg_fl_data_12_) );
	BUFX2 BUFX2_77 ( .A(data[13]), .Y(reg_fl_data_13_) );
	BUFX2 BUFX2_78 ( .A(data[14]), .Y(reg_fl_data_14_) );
	BUFX2 BUFX2_79 ( .A(data[15]), .Y(reg_fl_data_15_) );
	BUFX2 BUFX2_80 ( .A(clk), .Y(reg_fh_clk) );
	BUFX2 BUFX2_81 ( .A(reset), .Y(reg_fh_reset) );
	BUFX2 BUFX2_82 ( .A(data[0]), .Y(reg_vf_data_0_) );
	BUFX2 BUFX2_83 ( .A(data[1]), .Y(reg_vf_data_1_) );
	BUFX2 BUFX2_84 ( .A(data[2]), .Y(reg_vf_data_2_) );
	BUFX2 BUFX2_85 ( .A(data[3]), .Y(reg_vf_data_3_) );
	BUFX2 BUFX2_86 ( .A(data[4]), .Y(reg_vf_data_4_) );
	BUFX2 BUFX2_87 ( .A(data[5]), .Y(reg_vf_data_5_) );
	BUFX2 BUFX2_88 ( .A(data[6]), .Y(reg_vf_data_6_) );
	BUFX2 BUFX2_89 ( .A(data[7]), .Y(reg_vf_data_7_) );
	BUFX2 BUFX2_90 ( .A(data[8]), .Y(reg_vf_data_8_) );
	BUFX2 BUFX2_91 ( .A(data[9]), .Y(reg_vf_data_9_) );
	BUFX2 BUFX2_92 ( .A(data[10]), .Y(reg_vf_data_10_) );
	BUFX2 BUFX2_93 ( .A(data[11]), .Y(reg_vf_data_11_) );
	BUFX2 BUFX2_94 ( .A(data[12]), .Y(reg_vf_data_12_) );
	BUFX2 BUFX2_95 ( .A(data[13]), .Y(reg_vf_data_13_) );
	BUFX2 BUFX2_96 ( .A(data[14]), .Y(reg_vf_data_14_) );
	BUFX2 BUFX2_97 ( .A(data[15]), .Y(reg_vf_data_15_) );
	BUFX2 BUFX2_98 ( .A(addr_fh), .Y(reg_fh_cs) );
	BUFX2 BUFX2_99 ( .A(we), .Y(reg_fh_we) );
	BUFX2 BUFX2_100 ( .A(data[0]), .Y(reg_fh_data_0_) );
	BUFX2 BUFX2_101 ( .A(data[1]), .Y(reg_fh_data_1_) );
	BUFX2 BUFX2_102 ( .A(data[2]), .Y(reg_fh_data_2_) );
	BUFX2 BUFX2_103 ( .A(data[3]), .Y(reg_fh_data_3_) );
	BUFX2 BUFX2_104 ( .A(data[4]), .Y(reg_fh_data_4_) );
	BUFX2 BUFX2_105 ( .A(data[5]), .Y(reg_fh_data_5_) );
	BUFX2 BUFX2_106 ( .A(data[6]), .Y(reg_fh_data_6_) );
	BUFX2 BUFX2_107 ( .A(data[7]), .Y(reg_fh_data_7_) );
	BUFX2 BUFX2_108 ( .A(data[8]), .Y(reg_fh_data_8_) );
	BUFX2 BUFX2_109 ( .A(data[9]), .Y(reg_fh_data_9_) );
	BUFX2 BUFX2_110 ( .A(data[10]), .Y(reg_fh_data_10_) );
	BUFX2 BUFX2_111 ( .A(data[11]), .Y(reg_fh_data_11_) );
	BUFX2 BUFX2_112 ( .A(data[12]), .Y(reg_fh_data_12_) );
	BUFX2 BUFX2_113 ( .A(data[13]), .Y(reg_fh_data_13_) );
	BUFX2 BUFX2_114 ( .A(data[14]), .Y(reg_fh_data_14_) );
	BUFX2 BUFX2_115 ( .A(data[15]), .Y(reg_fh_data_15_) );
	BUFX2 BUFX2_116 ( .A(we), .Y(reg_vf_we) );
	BUFX2 BUFX2_117 ( .A(addr_vf), .Y(reg_vf_cs) );
	BUFX2 BUFX2_118 ( .A(reset), .Y(reg_vf_reset) );
	BUFX2 BUFX2_119 ( .A(clk), .Y(reg_vf_clk) );
	BUFX2 BUFX2_120 ( .A(data[0]), .Y(reg_ic_data_0_) );
	BUFX2 BUFX2_121 ( .A(data[1]), .Y(reg_ic_data_1_) );
	BUFX2 BUFX2_122 ( .A(data[2]), .Y(reg_ic_data_2_) );
	BUFX2 BUFX2_123 ( .A(data[3]), .Y(reg_ic_data_3_) );
	BUFX2 BUFX2_124 ( .A(data[4]), .Y(reg_ic_data_4_) );
	BUFX2 BUFX2_125 ( .A(data[5]), .Y(reg_ic_data_5_) );
	BUFX2 BUFX2_126 ( .A(data[6]), .Y(reg_ic_data_6_) );
	BUFX2 BUFX2_127 ( .A(data[7]), .Y(reg_ic_data_7_) );
	BUFX2 BUFX2_128 ( .A(data[8]), .Y(reg_ic_data_8_) );
	BUFX2 BUFX2_129 ( .A(data[9]), .Y(reg_ic_data_9_) );
	BUFX2 BUFX2_130 ( .A(data[10]), .Y(reg_ic_data_10_) );
	BUFX2 BUFX2_131 ( .A(data[11]), .Y(reg_ic_data_11_) );
	BUFX2 BUFX2_132 ( .A(data[12]), .Y(reg_ic_data_12_) );
	BUFX2 BUFX2_133 ( .A(data[13]), .Y(reg_ic_data_13_) );
	BUFX2 BUFX2_134 ( .A(data[14]), .Y(reg_ic_data_14_) );
	BUFX2 BUFX2_135 ( .A(data[15]), .Y(reg_ic_data_15_) );
	BUFX2 BUFX2_136 ( .A(we), .Y(reg_ic_we) );
	BUFX2 BUFX2_137 ( .A(addr_ic), .Y(reg_ic_cs) );
	BUFX2 BUFX2_138 ( .A(reset), .Y(reg_ic_reset) );
	BUFX2 BUFX2_139 ( .A(clk), .Y(reg_ic_clk) );
	BUFX2 BUFX2_140 ( .A(addr[0]), .Y(addr_decode_addr_0_) );
	BUFX2 BUFX2_141 ( .A(addr[1]), .Y(addr_decode_addr_1_) );
	BUFX2 BUFX2_142 ( .A(addr[2]), .Y(addr_decode_addr_2_) );
	BUFX2 BUFX2_143 ( .A(addr[3]), .Y(addr_decode_addr_3_) );
	BUFX2 BUFX2_144 ( .A(addr_hb), .Y(addr_decode_q_0_) );
	BUFX2 BUFX2_145 ( .A(addr_hv), .Y(addr_decode_q_1_) );
	BUFX2 BUFX2_146 ( .A(addr_hf), .Y(addr_decode_q_2_) );
	BUFX2 BUFX2_147 ( .A(addr_he), .Y(addr_decode_q_3_) );
	BUFX2 BUFX2_148 ( .A(addr_vb), .Y(addr_decode_q_4_) );
	BUFX2 BUFX2_149 ( .A(addr_vv), .Y(addr_decode_q_5_) );
	BUFX2 BUFX2_150 ( .A(addr_vf), .Y(addr_decode_q_6_) );
	BUFX2 BUFX2_151 ( .A(addr_ve), .Y(addr_decode_q_7_) );
	BUFX2 BUFX2_152 ( .A(addr_fl), .Y(addr_decode_q_8_) );
	BUFX2 BUFX2_153 ( .A(addr_fh), .Y(addr_decode_q_9_) );
	BUFX2 BUFX2_154 ( .A(addr_sl), .Y(addr_decode_q_10_) );
	BUFX2 BUFX2_155 ( .A(addr_sh), .Y(addr_decode_q_11_) );
	BUFX2 BUFX2_156 ( .A(addr_ic), .Y(addr_decode_q_12_) );
	BUFX2 BUFX2_157 ( .A(addr_ir), .Y(addr_decode_q_13_) );
	BUFX2 BUFX2_158 ( .A(addr_ia), .Y(addr_decode_q_14_) );
	BUFX2 BUFX2_159 ( .A(addr_cr), .Y(addr_decode_q_15_) );
	BUFX2 BUFX2_160 ( .A(data[0]), .Y(reg_vv_data_0_) );
	BUFX2 BUFX2_161 ( .A(data[1]), .Y(reg_vv_data_1_) );
	BUFX2 BUFX2_162 ( .A(data[2]), .Y(reg_vv_data_2_) );
	BUFX2 BUFX2_163 ( .A(data[3]), .Y(reg_vv_data_3_) );
	BUFX2 BUFX2_164 ( .A(data[4]), .Y(reg_vv_data_4_) );
	BUFX2 BUFX2_165 ( .A(data[5]), .Y(reg_vv_data_5_) );
	BUFX2 BUFX2_166 ( .A(data[6]), .Y(reg_vv_data_6_) );
	BUFX2 BUFX2_167 ( .A(data[7]), .Y(reg_vv_data_7_) );
	BUFX2 BUFX2_168 ( .A(data[8]), .Y(reg_vv_data_8_) );
	BUFX2 BUFX2_169 ( .A(data[9]), .Y(reg_vv_data_9_) );
	BUFX2 BUFX2_170 ( .A(data[10]), .Y(reg_vv_data_10_) );
	BUFX2 BUFX2_171 ( .A(data[11]), .Y(reg_vv_data_11_) );
	BUFX2 BUFX2_172 ( .A(data[12]), .Y(reg_vv_data_12_) );
	BUFX2 BUFX2_173 ( .A(data[13]), .Y(reg_vv_data_13_) );
	BUFX2 BUFX2_174 ( .A(data[14]), .Y(reg_vv_data_14_) );
	BUFX2 BUFX2_175 ( .A(data[15]), .Y(reg_vv_data_15_) );
	BUFX2 BUFX2_176 ( .A(we), .Y(reg_vv_we) );
	BUFX2 BUFX2_177 ( .A(addr_vv), .Y(reg_vv_cs) );
	BUFX2 BUFX2_178 ( .A(reset), .Y(reg_vv_reset) );
	BUFX2 BUFX2_179 ( .A(clk), .Y(reg_vv_clk) );
	BUFX2 BUFX2_180 ( .A(clk), .Y(reg_cr_clk) );
	BUFX2 BUFX2_181 ( .A(reset), .Y(reg_cr_reset) );
	BUFX2 BUFX2_182 ( .A(addr_cr), .Y(reg_cr_cs) );
	BUFX2 BUFX2_183 ( .A(we), .Y(reg_cr_we) );
	BUFX2 BUFX2_184 ( .A(data[0]), .Y(reg_cr_data_0_) );
	BUFX2 BUFX2_185 ( .A(data[1]), .Y(reg_cr_data_1_) );
	BUFX2 BUFX2_186 ( .A(data[2]), .Y(reg_cr_data_2_) );
	BUFX2 BUFX2_187 ( .A(data[3]), .Y(reg_cr_data_3_) );
	BUFX2 BUFX2_188 ( .A(data[4]), .Y(reg_cr_data_4_) );
	BUFX2 BUFX2_189 ( .A(data[5]), .Y(reg_cr_data_5_) );
	BUFX2 BUFX2_190 ( .A(data[6]), .Y(reg_cr_data_6_) );
	BUFX2 BUFX2_191 ( .A(data[7]), .Y(reg_cr_data_7_) );
	BUFX2 BUFX2_192 ( .A(data[8]), .Y(reg_cr_data_8_) );
	BUFX2 BUFX2_193 ( .A(data[9]), .Y(reg_cr_data_9_) );
	BUFX2 BUFX2_194 ( .A(data[10]), .Y(reg_cr_data_10_) );
	BUFX2 BUFX2_195 ( .A(data[11]), .Y(reg_cr_data_11_) );
	BUFX2 BUFX2_196 ( .A(data[12]), .Y(reg_cr_data_12_) );
	BUFX2 BUFX2_197 ( .A(data[13]), .Y(reg_cr_data_13_) );
	BUFX2 BUFX2_198 ( .A(data[14]), .Y(reg_cr_data_14_) );
	BUFX2 BUFX2_199 ( .A(data[15]), .Y(reg_cr_data_15_) );
	BUFX2 BUFX2_200 ( .A(data[0]), .Y(reg_vb_data_0_) );
	BUFX2 BUFX2_201 ( .A(data[1]), .Y(reg_vb_data_1_) );
	BUFX2 BUFX2_202 ( .A(data[2]), .Y(reg_vb_data_2_) );
	BUFX2 BUFX2_203 ( .A(data[3]), .Y(reg_vb_data_3_) );
	BUFX2 BUFX2_204 ( .A(data[4]), .Y(reg_vb_data_4_) );
	BUFX2 BUFX2_205 ( .A(data[5]), .Y(reg_vb_data_5_) );
	BUFX2 BUFX2_206 ( .A(data[6]), .Y(reg_vb_data_6_) );
	BUFX2 BUFX2_207 ( .A(data[7]), .Y(reg_vb_data_7_) );
	BUFX2 BUFX2_208 ( .A(data[8]), .Y(reg_vb_data_8_) );
	BUFX2 BUFX2_209 ( .A(data[9]), .Y(reg_vb_data_9_) );
	BUFX2 BUFX2_210 ( .A(data[10]), .Y(reg_vb_data_10_) );
	BUFX2 BUFX2_211 ( .A(data[11]), .Y(reg_vb_data_11_) );
	BUFX2 BUFX2_212 ( .A(data[12]), .Y(reg_vb_data_12_) );
	BUFX2 BUFX2_213 ( .A(data[13]), .Y(reg_vb_data_13_) );
	BUFX2 BUFX2_214 ( .A(data[14]), .Y(reg_vb_data_14_) );
	BUFX2 BUFX2_215 ( .A(data[15]), .Y(reg_vb_data_15_) );
	BUFX2 BUFX2_216 ( .A(we), .Y(reg_vb_we) );
	BUFX2 BUFX2_217 ( .A(addr_vb), .Y(reg_vb_cs) );
	BUFX2 BUFX2_218 ( .A(reset), .Y(reg_vb_reset) );
	BUFX2 BUFX2_219 ( .A(clk), .Y(reg_vb_clk) );
	BUFX2 BUFX2_220 ( .A(clk), .Y(reg_ir_clk) );
	BUFX2 BUFX2_221 ( .A(data[0]), .Y(reg_he_data_0_) );
	BUFX2 BUFX2_222 ( .A(data[1]), .Y(reg_he_data_1_) );
	BUFX2 BUFX2_223 ( .A(data[2]), .Y(reg_he_data_2_) );
	BUFX2 BUFX2_224 ( .A(data[3]), .Y(reg_he_data_3_) );
	BUFX2 BUFX2_225 ( .A(data[4]), .Y(reg_he_data_4_) );
	BUFX2 BUFX2_226 ( .A(data[5]), .Y(reg_he_data_5_) );
	BUFX2 BUFX2_227 ( .A(data[6]), .Y(reg_he_data_6_) );
	BUFX2 BUFX2_228 ( .A(data[7]), .Y(reg_he_data_7_) );
	BUFX2 BUFX2_229 ( .A(data[8]), .Y(reg_he_data_8_) );
	BUFX2 BUFX2_230 ( .A(data[9]), .Y(reg_he_data_9_) );
	BUFX2 BUFX2_231 ( .A(data[10]), .Y(reg_he_data_10_) );
	BUFX2 BUFX2_232 ( .A(data[11]), .Y(reg_he_data_11_) );
	BUFX2 BUFX2_233 ( .A(data[12]), .Y(reg_he_data_12_) );
	BUFX2 BUFX2_234 ( .A(data[13]), .Y(reg_he_data_13_) );
	BUFX2 BUFX2_235 ( .A(data[14]), .Y(reg_he_data_14_) );
	BUFX2 BUFX2_236 ( .A(data[15]), .Y(reg_he_data_15_) );
	BUFX2 BUFX2_237 ( .A(we), .Y(reg_he_we) );
	BUFX2 BUFX2_238 ( .A(addr_he), .Y(reg_he_cs) );
	BUFX2 BUFX2_239 ( .A(reset), .Y(reg_ir_reset) );
	BUFX2 BUFX2_240 ( .A(reset), .Y(reg_he_reset) );
	BUFX2 BUFX2_241 ( .A(clk), .Y(reg_he_clk) );
	BUFX2 BUFX2_242 ( .A(addr_ir), .Y(reg_ir_cs) );
	BUFX2 BUFX2_243 ( .A(we), .Y(reg_ir_we) );
	BUFX2 BUFX2_244 ( .A(clk), .Y(reg_sl_clk) );
	BUFX2 BUFX2_245 ( .A(reset), .Y(reg_sl_reset) );
	BUFX2 BUFX2_246 ( .A(addr_sl), .Y(reg_sl_cs) );
	BUFX2 BUFX2_247 ( .A(we), .Y(reg_sl_we) );
	BUFX2 BUFX2_248 ( .A(data[0]), .Y(reg_sl_data_0_) );
	BUFX2 BUFX2_249 ( .A(data[1]), .Y(reg_sl_data_1_) );
	BUFX2 BUFX2_250 ( .A(data[2]), .Y(reg_sl_data_2_) );
	BUFX2 BUFX2_251 ( .A(data[3]), .Y(reg_sl_data_3_) );
	BUFX2 BUFX2_252 ( .A(data[4]), .Y(reg_sl_data_4_) );
	BUFX2 BUFX2_253 ( .A(data[5]), .Y(reg_sl_data_5_) );
	BUFX2 BUFX2_254 ( .A(data[6]), .Y(reg_sl_data_6_) );
	BUFX2 BUFX2_255 ( .A(data[7]), .Y(reg_sl_data_7_) );
	BUFX2 BUFX2_256 ( .A(data[8]), .Y(reg_sl_data_8_) );
	BUFX2 BUFX2_257 ( .A(data[9]), .Y(reg_sl_data_9_) );
	BUFX2 BUFX2_258 ( .A(data[10]), .Y(reg_sl_data_10_) );
	BUFX2 BUFX2_259 ( .A(data[11]), .Y(reg_sl_data_11_) );
	BUFX2 BUFX2_260 ( .A(data[12]), .Y(reg_sl_data_12_) );
	BUFX2 BUFX2_261 ( .A(data[13]), .Y(reg_sl_data_13_) );
	BUFX2 BUFX2_262 ( .A(data[14]), .Y(reg_sl_data_14_) );
	BUFX2 BUFX2_263 ( .A(data[15]), .Y(reg_sl_data_15_) );
	BUFX2 BUFX2_264 ( .A(data[0]), .Y(reg_hf_data_0_) );
	BUFX2 BUFX2_265 ( .A(data[1]), .Y(reg_hf_data_1_) );
	BUFX2 BUFX2_266 ( .A(data[2]), .Y(reg_hf_data_2_) );
	BUFX2 BUFX2_267 ( .A(data[3]), .Y(reg_hf_data_3_) );
	BUFX2 BUFX2_268 ( .A(data[4]), .Y(reg_hf_data_4_) );
	BUFX2 BUFX2_269 ( .A(data[5]), .Y(reg_hf_data_5_) );
	BUFX2 BUFX2_270 ( .A(data[6]), .Y(reg_hf_data_6_) );
	BUFX2 BUFX2_271 ( .A(data[7]), .Y(reg_hf_data_7_) );
	BUFX2 BUFX2_272 ( .A(data[8]), .Y(reg_hf_data_8_) );
	BUFX2 BUFX2_273 ( .A(data[9]), .Y(reg_hf_data_9_) );
	BUFX2 BUFX2_274 ( .A(data[10]), .Y(reg_hf_data_10_) );
	BUFX2 BUFX2_275 ( .A(data[11]), .Y(reg_hf_data_11_) );
	BUFX2 BUFX2_276 ( .A(data[12]), .Y(reg_hf_data_12_) );
	BUFX2 BUFX2_277 ( .A(data[13]), .Y(reg_hf_data_13_) );
	BUFX2 BUFX2_278 ( .A(data[14]), .Y(reg_hf_data_14_) );
	BUFX2 BUFX2_279 ( .A(data[15]), .Y(reg_hf_data_15_) );
	BUFX2 BUFX2_280 ( .A(we), .Y(reg_hf_we) );
	BUFX2 BUFX2_281 ( .A(addr_hf), .Y(reg_hf_cs) );
	BUFX2 BUFX2_282 ( .A(reset), .Y(reg_hf_reset) );
	BUFX2 BUFX2_283 ( .A(clk), .Y(reg_hf_clk) );
	BUFX2 BUFX2_284 ( .A(data[0]), .Y(reg_hv_data_0_) );
	BUFX2 BUFX2_285 ( .A(data[1]), .Y(reg_hv_data_1_) );
	BUFX2 BUFX2_286 ( .A(data[2]), .Y(reg_hv_data_2_) );
	BUFX2 BUFX2_287 ( .A(data[3]), .Y(reg_hv_data_3_) );
	BUFX2 BUFX2_288 ( .A(data[4]), .Y(reg_hv_data_4_) );
	BUFX2 BUFX2_289 ( .A(data[5]), .Y(reg_hv_data_5_) );
	BUFX2 BUFX2_290 ( .A(data[6]), .Y(reg_hv_data_6_) );
	BUFX2 BUFX2_291 ( .A(data[7]), .Y(reg_hv_data_7_) );
	BUFX2 BUFX2_292 ( .A(data[8]), .Y(reg_hv_data_8_) );
	BUFX2 BUFX2_293 ( .A(data[9]), .Y(reg_hv_data_9_) );
	BUFX2 BUFX2_294 ( .A(data[10]), .Y(reg_hv_data_10_) );
	BUFX2 BUFX2_295 ( .A(data[11]), .Y(reg_hv_data_11_) );
	BUFX2 BUFX2_296 ( .A(data[12]), .Y(reg_hv_data_12_) );
	BUFX2 BUFX2_297 ( .A(data[13]), .Y(reg_hv_data_13_) );
	BUFX2 BUFX2_298 ( .A(data[14]), .Y(reg_hv_data_14_) );
	BUFX2 BUFX2_299 ( .A(data[15]), .Y(reg_hv_data_15_) );
	BUFX2 BUFX2_300 ( .A(we), .Y(reg_hv_we) );
	BUFX2 BUFX2_301 ( .A(addr_hv), .Y(reg_hv_cs) );
	BUFX2 BUFX2_302 ( .A(reset), .Y(reg_hv_reset) );
	BUFX2 BUFX2_303 ( .A(clk), .Y(reg_hv_clk) );
	BUFX2 BUFX2_304 ( .A(data[0]), .Y(reg_ir_data_0_) );
	BUFX2 BUFX2_305 ( .A(data[1]), .Y(reg_ir_data_1_) );
	BUFX2 BUFX2_306 ( .A(data[2]), .Y(reg_ir_data_2_) );
	BUFX2 BUFX2_307 ( .A(data[3]), .Y(reg_ir_data_3_) );
	BUFX2 BUFX2_308 ( .A(data[4]), .Y(reg_ir_data_4_) );
	BUFX2 BUFX2_309 ( .A(data[5]), .Y(reg_ir_data_5_) );
	BUFX2 BUFX2_310 ( .A(data[6]), .Y(reg_ir_data_6_) );
	BUFX2 BUFX2_311 ( .A(data[7]), .Y(reg_ir_data_7_) );
	BUFX2 BUFX2_312 ( .A(data[8]), .Y(reg_ir_data_8_) );
	BUFX2 BUFX2_313 ( .A(data[9]), .Y(reg_ir_data_9_) );
	BUFX2 BUFX2_314 ( .A(data[10]), .Y(reg_ir_data_10_) );
	BUFX2 BUFX2_315 ( .A(data[11]), .Y(reg_ir_data_11_) );
	BUFX2 BUFX2_316 ( .A(data[12]), .Y(reg_ir_data_12_) );
	BUFX2 BUFX2_317 ( .A(data[13]), .Y(reg_ir_data_13_) );
	BUFX2 BUFX2_318 ( .A(data[14]), .Y(reg_ir_data_14_) );
	BUFX2 BUFX2_319 ( .A(data[15]), .Y(reg_ir_data_15_) );
	BUFX2 BUFX2_320 ( .A(data[0]), .Y(reg_ve_data_0_) );
	BUFX2 BUFX2_321 ( .A(data[1]), .Y(reg_ve_data_1_) );
	BUFX2 BUFX2_322 ( .A(data[2]), .Y(reg_ve_data_2_) );
	BUFX2 BUFX2_323 ( .A(data[3]), .Y(reg_ve_data_3_) );
	BUFX2 BUFX2_324 ( .A(data[4]), .Y(reg_ve_data_4_) );
	BUFX2 BUFX2_325 ( .A(data[5]), .Y(reg_ve_data_5_) );
	BUFX2 BUFX2_326 ( .A(data[6]), .Y(reg_ve_data_6_) );
	BUFX2 BUFX2_327 ( .A(data[7]), .Y(reg_ve_data_7_) );
	BUFX2 BUFX2_328 ( .A(data[8]), .Y(reg_ve_data_8_) );
	BUFX2 BUFX2_329 ( .A(data[9]), .Y(reg_ve_data_9_) );
	BUFX2 BUFX2_330 ( .A(data[10]), .Y(reg_ve_data_10_) );
	BUFX2 BUFX2_331 ( .A(data[11]), .Y(reg_ve_data_11_) );
	BUFX2 BUFX2_332 ( .A(data[12]), .Y(reg_ve_data_12_) );
	BUFX2 BUFX2_333 ( .A(data[13]), .Y(reg_ve_data_13_) );
	BUFX2 BUFX2_334 ( .A(data[14]), .Y(reg_ve_data_14_) );
	BUFX2 BUFX2_335 ( .A(data[15]), .Y(reg_ve_data_15_) );
	BUFX2 BUFX2_336 ( .A(we), .Y(reg_ve_we) );
	BUFX2 BUFX2_337 ( .A(addr_ve), .Y(reg_ve_cs) );
	BUFX2 BUFX2_338 ( .A(reset), .Y(reg_ve_reset) );
	BUFX2 BUFX2_339 ( .A(clk), .Y(reg_ve_clk) );
	BUFX2 BUFX2_340 ( .A(reg_cr_value_5_), .Y(clk_select_0_) );
	BUFX2 BUFX2_341 ( .A(reg_cr_value_6_), .Y(clk_select_1_) );
	BUFX2 BUFX2_342 ( .A(reg_cr_value_7_), .Y(clk_select_2_) );
	BUFX2 BUFX2_343 ( .A(reg_cr_value_13_), .Y(vsync_invert) );
	BUFX2 BUFX2_344 ( .A(reg_cr_value_14_), .Y(hsync_invert) );
	BUFX2 BUFX2_345 ( .A(reg_cr_value_15_), .Y(irq_enabled) );
	BUFX2 BUFX2_346 ( .A(data[0]), .Y(reg_hb_data_0_) );
	BUFX2 BUFX2_347 ( .A(data[1]), .Y(reg_hb_data_1_) );
	BUFX2 BUFX2_348 ( .A(data[2]), .Y(reg_hb_data_2_) );
	BUFX2 BUFX2_349 ( .A(data[3]), .Y(reg_hb_data_3_) );
	BUFX2 BUFX2_350 ( .A(data[4]), .Y(reg_hb_data_4_) );
	BUFX2 BUFX2_351 ( .A(data[5]), .Y(reg_hb_data_5_) );
	BUFX2 BUFX2_352 ( .A(data[6]), .Y(reg_hb_data_6_) );
	BUFX2 BUFX2_353 ( .A(data[7]), .Y(reg_hb_data_7_) );
	BUFX2 BUFX2_354 ( .A(data[8]), .Y(reg_hb_data_8_) );
	BUFX2 BUFX2_355 ( .A(data[9]), .Y(reg_hb_data_9_) );
	BUFX2 BUFX2_356 ( .A(data[10]), .Y(reg_hb_data_10_) );
	BUFX2 BUFX2_357 ( .A(data[11]), .Y(reg_hb_data_11_) );
	BUFX2 BUFX2_358 ( .A(data[12]), .Y(reg_hb_data_12_) );
	BUFX2 BUFX2_359 ( .A(data[13]), .Y(reg_hb_data_13_) );
	BUFX2 BUFX2_360 ( .A(data[14]), .Y(reg_hb_data_14_) );
	BUFX2 BUFX2_361 ( .A(data[15]), .Y(reg_hb_data_15_) );
	BUFX2 BUFX2_362 ( .A(we), .Y(reg_hb_we) );
	BUFX2 BUFX2_363 ( .A(addr_hb), .Y(reg_hb_cs) );
	BUFX2 BUFX2_364 ( .A(reset), .Y(reg_hb_reset) );
	BUFX2 BUFX2_365 ( .A(reg_sl_value_0_), .Y(stride_0_) );
	BUFX2 BUFX2_366 ( .A(reg_sl_value_1_), .Y(stride_1_) );
	BUFX2 BUFX2_367 ( .A(reg_sl_value_2_), .Y(stride_2_) );
	BUFX2 BUFX2_368 ( .A(reg_sl_value_3_), .Y(stride_3_) );
	BUFX2 BUFX2_369 ( .A(reg_sl_value_4_), .Y(stride_4_) );
	BUFX2 BUFX2_370 ( .A(reg_sl_value_5_), .Y(stride_5_) );
	BUFX2 BUFX2_371 ( .A(reg_sl_value_6_), .Y(stride_6_) );
	BUFX2 BUFX2_372 ( .A(reg_sl_value_7_), .Y(stride_7_) );
	BUFX2 BUFX2_373 ( .A(reg_sl_value_8_), .Y(stride_8_) );
	BUFX2 BUFX2_374 ( .A(reg_sl_value_9_), .Y(stride_9_) );
	BUFX2 BUFX2_375 ( .A(reg_sl_value_10_), .Y(stride_10_) );
	BUFX2 BUFX2_376 ( .A(reg_sl_value_11_), .Y(stride_11_) );
	BUFX2 BUFX2_377 ( .A(reg_sl_value_12_), .Y(stride_12_) );
	BUFX2 BUFX2_378 ( .A(reg_sl_value_13_), .Y(stride_13_) );
	BUFX2 BUFX2_379 ( .A(reg_sl_value_14_), .Y(stride_14_) );
	BUFX2 BUFX2_380 ( .A(reg_sl_value_15_), .Y(stride_15_) );
	BUFX2 BUFX2_381 ( .A(reg_sh_value_0_), .Y(stride_16_) );
	BUFX2 BUFX2_382 ( .A(reg_sh_value_1_), .Y(stride_17_) );
	BUFX2 BUFX2_383 ( .A(reg_sh_value_2_), .Y(stride_18_) );
	BUFX2 BUFX2_384 ( .A(reg_sh_value_3_), .Y(stride_19_) );
	BUFX2 BUFX2_385 ( .A(reg_sh_value_4_), .Y(stride_20_) );
	BUFX2 BUFX2_386 ( .A(reg_sh_value_5_), .Y(stride_21_) );
	BUFX2 BUFX2_387 ( .A(reg_sh_value_6_), .Y(stride_22_) );
	BUFX2 BUFX2_388 ( .A(reg_sh_value_7_), .Y(stride_23_) );
	BUFX2 BUFX2_389 ( .A(reg_sh_value_8_), .Y(stride_24_) );
	BUFX2 BUFX2_390 ( .A(reg_sh_value_9_), .Y(stride_25_) );
	BUFX2 BUFX2_391 ( .A(reg_sh_value_10_), .Y(stride_26_) );
	BUFX2 BUFX2_392 ( .A(reg_sh_value_11_), .Y(stride_27_) );
	BUFX2 BUFX2_393 ( .A(reg_sh_value_12_), .Y(stride_28_) );
	BUFX2 BUFX2_394 ( .A(reg_sh_value_13_), .Y(stride_29_) );
	BUFX2 BUFX2_395 ( .A(reg_sh_value_14_), .Y(stride_30_) );
	BUFX2 BUFX2_396 ( .A(reg_sh_value_15_), .Y(stride_31_) );
	BUFX2 BUFX2_397 ( .A(reg_fl_value_0_), .Y(startaddr_0_) );
	BUFX2 BUFX2_398 ( .A(reg_fl_value_1_), .Y(startaddr_1_) );
	BUFX2 BUFX2_399 ( .A(reg_fl_value_2_), .Y(startaddr_2_) );
	BUFX2 BUFX2_400 ( .A(reg_fl_value_3_), .Y(startaddr_3_) );
	BUFX2 BUFX2_401 ( .A(reg_fl_value_4_), .Y(startaddr_4_) );
	BUFX2 BUFX2_402 ( .A(reg_fl_value_5_), .Y(startaddr_5_) );
	BUFX2 BUFX2_403 ( .A(reg_fl_value_6_), .Y(startaddr_6_) );
	BUFX2 BUFX2_404 ( .A(reg_fl_value_7_), .Y(startaddr_7_) );
	BUFX2 BUFX2_405 ( .A(reg_fl_value_8_), .Y(startaddr_8_) );
	BUFX2 BUFX2_406 ( .A(reg_fl_value_9_), .Y(startaddr_9_) );
	BUFX2 BUFX2_407 ( .A(reg_fl_value_10_), .Y(startaddr_10_) );
	BUFX2 BUFX2_408 ( .A(reg_fl_value_11_), .Y(startaddr_11_) );
	BUFX2 BUFX2_409 ( .A(reg_fl_value_12_), .Y(startaddr_12_) );
	BUFX2 BUFX2_410 ( .A(reg_fl_value_13_), .Y(startaddr_13_) );
	BUFX2 BUFX2_411 ( .A(reg_fl_value_14_), .Y(startaddr_14_) );
	BUFX2 BUFX2_412 ( .A(reg_fl_value_15_), .Y(startaddr_15_) );
	BUFX2 BUFX2_413 ( .A(reg_fh_value_0_), .Y(startaddr_16_) );
	BUFX2 BUFX2_414 ( .A(reg_fh_value_1_), .Y(startaddr_17_) );
	BUFX2 BUFX2_415 ( .A(reg_fh_value_2_), .Y(startaddr_18_) );
	BUFX2 BUFX2_416 ( .A(reg_fh_value_3_), .Y(startaddr_19_) );
	BUFX2 BUFX2_417 ( .A(reg_fh_value_4_), .Y(startaddr_20_) );
	BUFX2 BUFX2_418 ( .A(reg_fh_value_5_), .Y(startaddr_21_) );
	BUFX2 BUFX2_419 ( .A(reg_fh_value_6_), .Y(startaddr_22_) );
	BUFX2 BUFX2_420 ( .A(reg_fh_value_7_), .Y(startaddr_23_) );
	BUFX2 BUFX2_421 ( .A(reg_fh_value_8_), .Y(startaddr_24_) );
	BUFX2 BUFX2_422 ( .A(reg_fh_value_9_), .Y(startaddr_25_) );
	BUFX2 BUFX2_423 ( .A(reg_fh_value_10_), .Y(startaddr_26_) );
	BUFX2 BUFX2_424 ( .A(reg_fh_value_11_), .Y(startaddr_27_) );
	BUFX2 BUFX2_425 ( .A(reg_fh_value_12_), .Y(startaddr_28_) );
	BUFX2 BUFX2_426 ( .A(reg_fh_value_13_), .Y(startaddr_29_) );
	BUFX2 BUFX2_427 ( .A(reg_fh_value_14_), .Y(startaddr_30_) );
	BUFX2 BUFX2_428 ( .A(reg_fh_value_15_), .Y(startaddr_31_) );
	BUFX2 BUFX2_429 ( .A(reg_cr_value_0_), .Y(control_0_) );
	BUFX2 BUFX2_430 ( .A(reg_cr_value_1_), .Y(control_1_) );
	BUFX2 BUFX2_431 ( .A(reg_cr_value_2_), .Y(control_2_) );
	BUFX2 BUFX2_432 ( .A(reg_cr_value_3_), .Y(control_3_) );
	BUFX2 BUFX2_433 ( .A(reg_cr_value_4_), .Y(control_4_) );
	BUFX2 BUFX2_434 ( .A(reg_cr_value_5_), .Y(control_5_) );
	BUFX2 BUFX2_435 ( .A(reg_cr_value_6_), .Y(control_6_) );
	BUFX2 BUFX2_436 ( .A(reg_cr_value_7_), .Y(control_7_) );
	BUFX2 BUFX2_437 ( .A(reg_cr_value_8_), .Y(control_8_) );
	BUFX2 BUFX2_438 ( .A(reg_cr_value_9_), .Y(control_9_) );
	BUFX2 BUFX2_439 ( .A(reg_cr_value_10_), .Y(control_10_) );
	BUFX2 BUFX2_440 ( .A(reg_cr_value_11_), .Y(control_11_) );
	BUFX2 BUFX2_441 ( .A(reg_cr_value_12_), .Y(control_12_) );
	BUFX2 BUFX2_442 ( .A(reg_cr_value_13_), .Y(control_13_) );
	BUFX2 BUFX2_443 ( .A(reg_cr_value_14_), .Y(control_14_) );
	BUFX2 BUFX2_444 ( .A(reg_cr_value_15_), .Y(control_15_) );
	BUFX2 BUFX2_445 ( .A(reg_ir_value_0_), .Y(irqr_0_) );
	BUFX2 BUFX2_446 ( .A(reg_ir_value_1_), .Y(irqr_1_) );
	BUFX2 BUFX2_447 ( .A(reg_ir_value_2_), .Y(irqr_2_) );
	BUFX2 BUFX2_448 ( .A(reg_ir_value_3_), .Y(irqr_3_) );
	BUFX2 BUFX2_449 ( .A(reg_ir_value_4_), .Y(irqr_4_) );
	BUFX2 BUFX2_450 ( .A(reg_ir_value_5_), .Y(irqr_5_) );
	BUFX2 BUFX2_451 ( .A(reg_ir_value_6_), .Y(irqr_6_) );
	BUFX2 BUFX2_452 ( .A(reg_ir_value_7_), .Y(irqr_7_) );
	BUFX2 BUFX2_453 ( .A(reg_ir_value_8_), .Y(irqr_8_) );
	BUFX2 BUFX2_454 ( .A(reg_ir_value_9_), .Y(irqr_9_) );
	BUFX2 BUFX2_455 ( .A(reg_ir_value_10_), .Y(irqr_10_) );
	BUFX2 BUFX2_456 ( .A(reg_ir_value_11_), .Y(irqr_11_) );
	BUFX2 BUFX2_457 ( .A(reg_ir_value_12_), .Y(irqr_12_) );
	BUFX2 BUFX2_458 ( .A(reg_ir_value_13_), .Y(irqr_13_) );
	BUFX2 BUFX2_459 ( .A(reg_ir_value_14_), .Y(irqr_14_) );
	BUFX2 BUFX2_460 ( .A(reg_ir_value_15_), .Y(irqr_15_) );
	BUFX2 BUFX2_461 ( .A(reg_ic_value_0_), .Y(irqc_0_) );
	BUFX2 BUFX2_462 ( .A(reg_ic_value_1_), .Y(irqc_1_) );
	BUFX2 BUFX2_463 ( .A(reg_ic_value_2_), .Y(irqc_2_) );
	BUFX2 BUFX2_464 ( .A(reg_ic_value_3_), .Y(irqc_3_) );
	BUFX2 BUFX2_465 ( .A(reg_ic_value_4_), .Y(irqc_4_) );
	BUFX2 BUFX2_466 ( .A(reg_ic_value_5_), .Y(irqc_5_) );
	BUFX2 BUFX2_467 ( .A(reg_ic_value_6_), .Y(irqc_6_) );
	BUFX2 BUFX2_468 ( .A(reg_ic_value_7_), .Y(irqc_7_) );
	BUFX2 BUFX2_469 ( .A(reg_ic_value_8_), .Y(irqc_8_) );
	BUFX2 BUFX2_470 ( .A(reg_ic_value_9_), .Y(irqc_9_) );
	BUFX2 BUFX2_471 ( .A(reg_ic_value_10_), .Y(irqc_10_) );
	BUFX2 BUFX2_472 ( .A(reg_ic_value_11_), .Y(irqc_11_) );
	BUFX2 BUFX2_473 ( .A(reg_ic_value_12_), .Y(irqc_12_) );
	BUFX2 BUFX2_474 ( .A(reg_ic_value_13_), .Y(irqc_13_) );
	BUFX2 BUFX2_475 ( .A(reg_ic_value_14_), .Y(irqc_14_) );
	BUFX2 BUFX2_476 ( .A(reg_ic_value_15_), .Y(irqc_15_) );
	BUFX2 BUFX2_477 ( .A(reg_ve_value_0_), .Y(vend_0_) );
	BUFX2 BUFX2_478 ( .A(reg_ve_value_1_), .Y(vend_1_) );
	BUFX2 BUFX2_479 ( .A(reg_ve_value_2_), .Y(vend_2_) );
	BUFX2 BUFX2_480 ( .A(reg_ve_value_3_), .Y(vend_3_) );
	BUFX2 BUFX2_481 ( .A(reg_ve_value_4_), .Y(vend_4_) );
	BUFX2 BUFX2_482 ( .A(reg_ve_value_5_), .Y(vend_5_) );
	BUFX2 BUFX2_483 ( .A(reg_ve_value_6_), .Y(vend_6_) );
	BUFX2 BUFX2_484 ( .A(reg_ve_value_7_), .Y(vend_7_) );
	BUFX2 BUFX2_485 ( .A(reg_ve_value_8_), .Y(vend_8_) );
	BUFX2 BUFX2_486 ( .A(reg_ve_value_9_), .Y(vend_9_) );
	BUFX2 BUFX2_487 ( .A(reg_ve_value_10_), .Y(vend_10_) );
	BUFX2 BUFX2_488 ( .A(reg_ve_value_11_), .Y(vend_11_) );
	BUFX2 BUFX2_489 ( .A(reg_ve_value_12_), .Y(vend_12_) );
	BUFX2 BUFX2_490 ( .A(reg_ve_value_13_), .Y(vend_13_) );
	BUFX2 BUFX2_491 ( .A(reg_ve_value_14_), .Y(vend_14_) );
	BUFX2 BUFX2_492 ( .A(reg_ve_value_15_), .Y(vend_15_) );
	BUFX2 BUFX2_493 ( .A(reg_vf_value_0_), .Y(vfporch_0_) );
	BUFX2 BUFX2_494 ( .A(reg_vf_value_1_), .Y(vfporch_1_) );
	BUFX2 BUFX2_495 ( .A(reg_vf_value_2_), .Y(vfporch_2_) );
	BUFX2 BUFX2_496 ( .A(reg_vf_value_3_), .Y(vfporch_3_) );
	BUFX2 BUFX2_497 ( .A(reg_vf_value_4_), .Y(vfporch_4_) );
	BUFX2 BUFX2_498 ( .A(reg_vf_value_5_), .Y(vfporch_5_) );
	BUFX2 BUFX2_499 ( .A(reg_vf_value_6_), .Y(vfporch_6_) );
	BUFX2 BUFX2_500 ( .A(reg_vf_value_7_), .Y(vfporch_7_) );
	BUFX2 BUFX2_501 ( .A(reg_vf_value_8_), .Y(vfporch_8_) );
	BUFX2 BUFX2_502 ( .A(reg_vf_value_9_), .Y(vfporch_9_) );
	BUFX2 BUFX2_503 ( .A(reg_vf_value_10_), .Y(vfporch_10_) );
	BUFX2 BUFX2_504 ( .A(reg_vf_value_11_), .Y(vfporch_11_) );
	BUFX2 BUFX2_505 ( .A(reg_vf_value_12_), .Y(vfporch_12_) );
	BUFX2 BUFX2_506 ( .A(reg_vf_value_13_), .Y(vfporch_13_) );
	BUFX2 BUFX2_507 ( .A(reg_vf_value_14_), .Y(vfporch_14_) );
	BUFX2 BUFX2_508 ( .A(reg_vf_value_15_), .Y(vfporch_15_) );
	BUFX2 BUFX2_509 ( .A(reg_vv_value_0_), .Y(vvideo_0_) );
	BUFX2 BUFX2_510 ( .A(reg_vv_value_1_), .Y(vvideo_1_) );
	BUFX2 BUFX2_511 ( .A(reg_vv_value_2_), .Y(vvideo_2_) );
	BUFX2 BUFX2_512 ( .A(reg_vv_value_3_), .Y(vvideo_3_) );
	BUFX2 BUFX2_513 ( .A(reg_vv_value_4_), .Y(vvideo_4_) );
	BUFX2 BUFX2_514 ( .A(reg_vv_value_5_), .Y(vvideo_5_) );
	BUFX2 BUFX2_515 ( .A(reg_vv_value_6_), .Y(vvideo_6_) );
	BUFX2 BUFX2_516 ( .A(reg_vv_value_7_), .Y(vvideo_7_) );
	BUFX2 BUFX2_517 ( .A(reg_vv_value_8_), .Y(vvideo_8_) );
	BUFX2 BUFX2_518 ( .A(reg_vv_value_9_), .Y(vvideo_9_) );
	BUFX2 BUFX2_519 ( .A(reg_vv_value_10_), .Y(vvideo_10_) );
	BUFX2 BUFX2_520 ( .A(reg_vv_value_11_), .Y(vvideo_11_) );
	BUFX2 BUFX2_521 ( .A(reg_vv_value_12_), .Y(vvideo_12_) );
	BUFX2 BUFX2_522 ( .A(reg_vv_value_13_), .Y(vvideo_13_) );
	BUFX2 BUFX2_523 ( .A(reg_vv_value_14_), .Y(vvideo_14_) );
	BUFX2 BUFX2_524 ( .A(reg_vv_value_15_), .Y(vvideo_15_) );
	BUFX2 BUFX2_525 ( .A(reg_vb_value_0_), .Y(vbporch_0_) );
	BUFX2 BUFX2_526 ( .A(reg_vb_value_1_), .Y(vbporch_1_) );
	BUFX2 BUFX2_527 ( .A(reg_vb_value_2_), .Y(vbporch_2_) );
	BUFX2 BUFX2_528 ( .A(reg_vb_value_3_), .Y(vbporch_3_) );
	BUFX2 BUFX2_529 ( .A(reg_vb_value_4_), .Y(vbporch_4_) );
	BUFX2 BUFX2_530 ( .A(reg_vb_value_5_), .Y(vbporch_5_) );
	BUFX2 BUFX2_531 ( .A(reg_vb_value_6_), .Y(vbporch_6_) );
	BUFX2 BUFX2_532 ( .A(reg_vb_value_7_), .Y(vbporch_7_) );
	BUFX2 BUFX2_533 ( .A(reg_vb_value_8_), .Y(vbporch_8_) );
	BUFX2 BUFX2_534 ( .A(reg_vb_value_9_), .Y(vbporch_9_) );
	BUFX2 BUFX2_535 ( .A(reg_vb_value_10_), .Y(vbporch_10_) );
	BUFX2 BUFX2_536 ( .A(reg_vb_value_11_), .Y(vbporch_11_) );
	BUFX2 BUFX2_537 ( .A(reg_vb_value_12_), .Y(vbporch_12_) );
	BUFX2 BUFX2_538 ( .A(reg_vb_value_13_), .Y(vbporch_13_) );
	BUFX2 BUFX2_539 ( .A(reg_vb_value_14_), .Y(vbporch_14_) );
	BUFX2 BUFX2_540 ( .A(reg_vb_value_15_), .Y(vbporch_15_) );
	BUFX2 BUFX2_541 ( .A(reg_he_value_0_), .Y(hend_0_) );
	BUFX2 BUFX2_542 ( .A(reg_he_value_1_), .Y(hend_1_) );
	BUFX2 BUFX2_543 ( .A(reg_he_value_2_), .Y(hend_2_) );
	BUFX2 BUFX2_544 ( .A(reg_he_value_3_), .Y(hend_3_) );
	BUFX2 BUFX2_545 ( .A(reg_he_value_4_), .Y(hend_4_) );
	BUFX2 BUFX2_546 ( .A(reg_he_value_5_), .Y(hend_5_) );
	BUFX2 BUFX2_547 ( .A(reg_he_value_6_), .Y(hend_6_) );
	BUFX2 BUFX2_548 ( .A(reg_he_value_7_), .Y(hend_7_) );
	BUFX2 BUFX2_549 ( .A(reg_he_value_8_), .Y(hend_8_) );
	BUFX2 BUFX2_550 ( .A(reg_he_value_9_), .Y(hend_9_) );
	BUFX2 BUFX2_551 ( .A(reg_he_value_10_), .Y(hend_10_) );
	BUFX2 BUFX2_552 ( .A(reg_he_value_11_), .Y(hend_11_) );
	BUFX2 BUFX2_553 ( .A(reg_he_value_12_), .Y(hend_12_) );
	BUFX2 BUFX2_554 ( .A(reg_he_value_13_), .Y(hend_13_) );
	BUFX2 BUFX2_555 ( .A(reg_he_value_14_), .Y(hend_14_) );
	BUFX2 BUFX2_556 ( .A(reg_he_value_15_), .Y(hend_15_) );
	BUFX2 BUFX2_557 ( .A(reg_hf_value_0_), .Y(hfporch_0_) );
	BUFX2 BUFX2_558 ( .A(reg_hf_value_1_), .Y(hfporch_1_) );
	BUFX2 BUFX2_559 ( .A(reg_hf_value_2_), .Y(hfporch_2_) );
	BUFX2 BUFX2_560 ( .A(reg_hf_value_3_), .Y(hfporch_3_) );
	BUFX2 BUFX2_561 ( .A(reg_hf_value_4_), .Y(hfporch_4_) );
	BUFX2 BUFX2_562 ( .A(reg_hf_value_5_), .Y(hfporch_5_) );
	BUFX2 BUFX2_563 ( .A(reg_hf_value_6_), .Y(hfporch_6_) );
	BUFX2 BUFX2_564 ( .A(reg_hf_value_7_), .Y(hfporch_7_) );
	BUFX2 BUFX2_565 ( .A(reg_hf_value_8_), .Y(hfporch_8_) );
	BUFX2 BUFX2_566 ( .A(reg_hf_value_9_), .Y(hfporch_9_) );
	BUFX2 BUFX2_567 ( .A(reg_hf_value_10_), .Y(hfporch_10_) );
	BUFX2 BUFX2_568 ( .A(reg_hf_value_11_), .Y(hfporch_11_) );
	BUFX2 BUFX2_569 ( .A(reg_hf_value_12_), .Y(hfporch_12_) );
	BUFX2 BUFX2_570 ( .A(reg_hf_value_13_), .Y(hfporch_13_) );
	BUFX2 BUFX2_571 ( .A(reg_hf_value_14_), .Y(hfporch_14_) );
	BUFX2 BUFX2_572 ( .A(reg_hf_value_15_), .Y(hfporch_15_) );
	BUFX2 BUFX2_573 ( .A(reg_hv_value_0_), .Y(hvideo_0_) );
	BUFX2 BUFX2_574 ( .A(reg_hv_value_1_), .Y(hvideo_1_) );
	BUFX2 BUFX2_575 ( .A(reg_hv_value_2_), .Y(hvideo_2_) );
	BUFX2 BUFX2_576 ( .A(reg_hv_value_3_), .Y(hvideo_3_) );
	BUFX2 BUFX2_577 ( .A(reg_hv_value_4_), .Y(hvideo_4_) );
	BUFX2 BUFX2_578 ( .A(reg_hv_value_5_), .Y(hvideo_5_) );
	BUFX2 BUFX2_579 ( .A(reg_hv_value_6_), .Y(hvideo_6_) );
	BUFX2 BUFX2_580 ( .A(reg_hv_value_7_), .Y(hvideo_7_) );
	BUFX2 BUFX2_581 ( .A(reg_hv_value_8_), .Y(hvideo_8_) );
	BUFX2 BUFX2_582 ( .A(reg_hv_value_9_), .Y(hvideo_9_) );
	BUFX2 BUFX2_583 ( .A(reg_hv_value_10_), .Y(hvideo_10_) );
	BUFX2 BUFX2_584 ( .A(reg_hv_value_11_), .Y(hvideo_11_) );
	BUFX2 BUFX2_585 ( .A(reg_hv_value_12_), .Y(hvideo_12_) );
	BUFX2 BUFX2_586 ( .A(reg_hv_value_13_), .Y(hvideo_13_) );
	BUFX2 BUFX2_587 ( .A(reg_hv_value_14_), .Y(hvideo_14_) );
	BUFX2 BUFX2_588 ( .A(reg_hv_value_15_), .Y(hvideo_15_) );
	BUFX2 BUFX2_589 ( .A(reg_hb_value_0_), .Y(hbporch_0_) );
	BUFX2 BUFX2_590 ( .A(reg_hb_value_1_), .Y(hbporch_1_) );
	BUFX2 BUFX2_591 ( .A(reg_hb_value_2_), .Y(hbporch_2_) );
	BUFX2 BUFX2_592 ( .A(reg_hb_value_3_), .Y(hbporch_3_) );
	BUFX2 BUFX2_593 ( .A(reg_hb_value_4_), .Y(hbporch_4_) );
	BUFX2 BUFX2_594 ( .A(reg_hb_value_5_), .Y(hbporch_5_) );
	BUFX2 BUFX2_595 ( .A(reg_hb_value_6_), .Y(hbporch_6_) );
	BUFX2 BUFX2_596 ( .A(reg_hb_value_7_), .Y(hbporch_7_) );
	BUFX2 BUFX2_597 ( .A(reg_hb_value_8_), .Y(hbporch_8_) );
	BUFX2 BUFX2_598 ( .A(reg_hb_value_9_), .Y(hbporch_9_) );
	BUFX2 BUFX2_599 ( .A(reg_hb_value_10_), .Y(hbporch_10_) );
	BUFX2 BUFX2_600 ( .A(reg_hb_value_11_), .Y(hbporch_11_) );
	BUFX2 BUFX2_601 ( .A(reg_hb_value_12_), .Y(hbporch_12_) );
	BUFX2 BUFX2_602 ( .A(reg_hb_value_13_), .Y(hbporch_13_) );
	BUFX2 BUFX2_603 ( .A(reg_hb_value_14_), .Y(hbporch_14_) );
	BUFX2 BUFX2_604 ( .A(reg_hb_value_15_), .Y(hbporch_15_) );
	BUFX2 BUFX2_605 ( .A(clk), .Y(reg_hb_clk) );
endmodule
